32'sd191286, 32'sd363208, 32'sd350652, 32'sd504747, 32'sd398543, 32'sd210904, 32'sd277821, 32'sd177590, 32'sd878147, 32'sd333487,
32'sd5678, 32'sd338304, 32'sd106838, 32'sd9669, 32'sd437062, 32'sd918260, 32'sd215831, 32'sd114457, 32'sd231213, 32'sd83398,
32'sd144142, 32'sd337134, 32'sd549572, 32'sd501385, 32'sd16821, 32'sd229739, 32'sd7410, 32'sd132301, 32'sd311534, 32'sd238326,
32'sd107294, 32'sd57729, 32'sd20423, 32'sd140663, 32'sd228067, 32'sd104717, 32'sd448416, 32'sd266303, 32'sd964782, 32'sd351866,
32'sd558936, 32'sd505616, 32'sd173238, 32'sd181845, 32'sd159025, 32'sd359747, 32'sd191896, 32'sd414635, 32'sd44897, 32'sd3346,
32'sd257100, 32'sd210885, 32'sd66293, 32'sd63400, 32'sd189979, 32'sd77144, 32'sd163564, 32'sd599407, 32'sd668735, 32'sd216124,
32'sd87853, 32'sd302209, 32'sd493297, 32'sd331451, 32'sd35441, 32'sd270547, 32'sd248656, 32'sd443469, 32'sd45373, 32'sd378831,
32'sd509375, 32'sd227772, 32'sd21172, 32'sd16396, 32'sd194124, 32'sd4273, 32'sd24766, 32'sd579178, 32'sd115658, 32'sd74515,
32'sd19350, 32'sd148397, 32'sd179174, 32'sd90723, 32'sd57463, 32'sd451867, 32'sd256552, 32'sd161100, 32'sd756940, 32'sd477810,
32'sd78573, 32'sd21474, 32'sd189698, 32'sd422517, 32'sd66385, 32'sd295243, 32'sd345735, 32'sd133455, 32'sd62002, 32'sd143020,
32'sd334033, 32'sd227439, 32'sd691911, 32'sd339279, 32'sd102660, 32'sd511061, 32'sd611219, 32'sd796154, 32'sd198799, 32'sd77415,
32'sd17150, 32'sd221695, 32'sd57099, 32'sd464501, 32'sd341712, 32'sd186041, 32'sd25343, 32'sd202833, 32'sd122656, 32'sd297849,
32'sd465216, 32'sd44400, 32'sd854290, 32'sd47654, 32'sd790356, 32'sd285316, 32'sd672401, 32'sd74602, 32'sd108750, 32'sd55939,
32'sd101380, 32'sd244424, 32'sd236, 32'sd488225, 32'sd195103, 32'sd199795, 32'sd191447, 32'sd201105, 32'sd352346, 32'sd37528,
32'sd478545, 32'sd469462, 32'sd605691, 32'sd162573, 32'sd478763, 32'sd85437, 32'sd69509, 32'sd111452, 32'sd138211, 32'sd363984,
32'sd149779, 32'sd149864, 32'sd557572, 32'sd4136, 32'sd898730, 32'sd309180, 32'sd143859, 32'sd211501, 32'sd158090, 32'sd186506,
32'sd216647, 32'sd314787, 32'sd337857, 32'sd392551, 32'sd156862, 32'sd487599, 32'sd46665, 32'sd345355, 32'sd269421, 32'sd89943,
32'sd492773, 32'sd888818, 32'sd60794, 32'sd288313, 32'sd646823, 32'sd131297, 32'sd447130, 32'sd472611, 32'sd234237, 32'sd63906,
32'sd1096984, 32'sd494849, 32'sd146363, 32'sd4214, 32'sd399348, 32'sd108992, 32'sd26001, 32'sd312840, 32'sd60253, 32'sd268636,
32'sd365674, 32'sd75835, 32'sd449673, 32'sd3322, 32'sd589784, 32'sd379912, 32'sd388146, 32'sd149765, 32'sd15694, 32'sd538533,
32'sd130963, 32'sd919122, 32'sd5397, 32'sd46922, 32'sd544932, 32'sd413191, 32'sd185923, 32'sd27043, 32'sd46667, 32'sd634659,
32'sd795075, 32'sd102362, 32'sd19705, 32'sd812497, 32'sd259981, 32'sd1384694, 32'sd31353, 32'sd196933, 32'sd186321, 32'sd314916,
32'sd14363, 32'sd106245, 32'sd111345, 32'sd34711, 32'sd56854, 32'sd20679, 32'sd459078, 32'sd110582, 32'sd41448, 32'sd66571,
32'sd666064, 32'sd765109, 32'sd141930, 32'sd144157, 32'sd41724, 32'sd8435, 32'sd26856, 32'sd44489, 32'sd95625, 32'sd663275,
32'sd1098622, 32'sd524796, 32'sd342016, 32'sd1069536, 32'sd277828, 32'sd311159, 32'sd370749, 32'sd479785, 32'sd241792, 32'sd476030,
32'sd1356964, 32'sd28527, 32'sd301825, 32'sd219837, 32'sd51442, 32'sd159882, 32'sd130956, 32'sd50102, 32'sd248481, 32'sd53532,
32'sd510823, 32'sd95798, 32'sd785289, 32'sd159975, 32'sd74293, 32'sd314985, 32'sd255958, 32'sd240449, 32'sd698015, 32'sd671580,
32'sd116794, 32'sd142964, 32'sd99378, 32'sd251040, 32'sd55434, 32'sd558858, 32'sd270148, 32'sd22786, 32'sd157852, 32'sd245697,
32'sd48541, 32'sd133851, 32'sd357273, 32'sd242102, 32'sd133085, 32'sd340023, 32'sd175634, 32'sd216452, 32'sd9449, 32'sd496786,
32'sd425419, 32'sd166801, 32'sd88543, 32'sd241363, 32'sd227444, 32'sd34976, 32'sd246468, 32'sd70474, 32'sd57609, 32'sd41473,
32'sd660346, 32'sd466905, 32'sd159846, 32'sd694368, 32'sd459816, 32'sd77950, 32'sd234785, 32'sd292897, 32'sd294944, 32'sd568667,
32'sd407242, 32'sd1013895, 32'sd357045, 32'sd61320, 32'sd218197, 32'sd206602, 32'sd137624, 32'sd110752, 32'sd73440, 32'sd111768,
32'sd473920, 32'sd161456, 32'sd125590, 32'sd562068, 32'sd238180, 32'sd298383, 32'sd225699, 32'sd274029, 32'sd648883, 32'sd201831,
32'sd163891, 32'sd265537, 32'sd324881, 32'sd74425, 32'sd210260, 32'sd118736, 32'sd381134, 32'sd129400, 32'sd405163, 32'sd22616,
32'sd129035, 32'sd319443, 32'sd98203, 32'sd848882, 32'sd76061, 32'sd242786, 32'sd163611, 32'sd451526, 32'sd28604, 32'sd408109,
32'sd843115, 32'sd32642, 32'sd362070, 32'sd372841, 32'sd196056, 32'sd364105, 32'sd272173, 32'sd410421, 32'sd737722, 32'sd219316,
32'sd237101, 32'sd97720, 32'sd309434, 32'sd283316, 32'sd392480, 32'sd22050, 32'sd228688, 32'sd140496, 32'sd61548, 32'sd291123,
32'sd304398, 32'sd331439, 32'sd252151, 32'sd66943, 32'sd69414, 32'sd234259, 32'sd569479, 32'sd22698, 32'sd77227, 32'sd263261,
32'sd140482, 32'sd126717, 32'sd501925, 32'sd239386, 32'sd169253, 32'sd2453, 32'sd125268, 32'sd39587, 32'sd230930, 32'sd275010,
32'sd119618, 32'sd253603, 32'sd329629, 32'sd831427, 32'sd202578, 32'sd365900, 32'sd311423, 32'sd493272, 32'sd594497, 32'sd132279,
32'sd89617, 32'sd266151, 32'sd58217, 32'sd645832, 32'sd476502, 32'sd312456, 32'sd33487, 32'sd17189, 32'sd69097, 32'sd407085,
32'sd222260, 32'sd125279, 32'sd57252, 32'sd683692, 32'sd100461, 32'sd148998, 32'sd262178, 32'sd120143, 32'sd13242, 32'sd235544,
32'sd123927, 32'sd5803, 32'sd154176, 32'sd421486, 32'sd416630, 32'sd7647, 32'sd219182, 32'sd405981, 32'sd390648, 32'sd12127,
32'sd8422, 32'sd370018, 32'sd660488, 32'sd164410, 32'sd181835, 32'sd170600, 32'sd304834, 32'sd149593, 32'sd520128, 32'sd131054,
32'sd139513, 32'sd652881, 32'sd242039, 32'sd767896, 32'sd523267, 32'sd388355, 32'sd411593, 32'sd300627, 32'sd770185, 32'sd621289,
32'sd189727, 32'sd144564, 32'sd80442, 32'sd150537, 32'sd277756, 32'sd679687, 32'sd646952, 32'sd190922, 32'sd19597, 32'sd67521,
32'sd271146, 32'sd224144, 32'sd263508, 32'sd240668, 32'sd102517, 32'sd609665, 32'sd208983, 32'sd565127, 32'sd462249, 32'sd218046,
32'sd17440, 32'sd582208, 32'sd170686, 32'sd4277, 32'sd193569, 32'sd176692, 32'sd361080, 32'sd24403, 32'sd235851, 32'sd594113,
32'sd27298, 32'sd110237, 32'sd26663, 32'sd308360, 32'sd582469, 32'sd560986, 32'sd359285, 32'sd311309, 32'sd207163, 32'sd33073,
32'sd36226, 32'sd128421, 32'sd153882, 32'sd111492, 32'sd84902, 32'sd470213, 32'sd842329, 32'sd292793, 32'sd52963, 32'sd139279,
32'sd242335, 32'sd129037, 32'sd29079, 32'sd105655, 32'sd149888, 32'sd516363, 32'sd740994, 32'sd207092, 32'sd161196, 32'sd156753,
32'sd315808, 32'sd673194, 32'sd141604, 32'sd752182, 32'sd795893, 32'sd197472, 32'sd130730, 32'sd64603, 32'sd991174, 32'sd82479,
32'sd213604, 32'sd647257, 32'sd701810, 32'sd368060, 32'sd201463, 32'sd207751, 32'sd140040, 32'sd196701, 32'sd394050, 32'sd112758,
32'sd152347, 32'sd499457, 32'sd160915, 32'sd89698, 32'sd171124, 32'sd48213, 32'sd295109, 32'sd173961, 32'sd1028340, 32'sd432796,
32'sd8910, 32'sd401324, 32'sd122398, 32'sd580058, 32'sd75363, 32'sd280236, 32'sd6860, 32'sd51475, 32'sd827054, 32'sd366968,
32'sd562089, 32'sd431780, 32'sd89663, 32'sd317330, 32'sd2149, 32'sd236430, 32'sd141370, 32'sd32645, 32'sd130886, 32'sd426441,
32'sd97896, 32'sd91983, 32'sd133318, 32'sd2732, 32'sd133598, 32'sd1235650, 32'sd378148, 32'sd180202, 32'sd55973, 32'sd388115,
32'sd57968, 32'sd288499, 32'sd113120, 32'sd83528, 32'sd154895, 32'sd40920, 32'sd153423, 32'sd26541, 32'sd162801, 32'sd148736,
32'sd34357, 32'sd305791, 32'sd580369, 32'sd141150, 32'sd82144, 32'sd86448, 32'sd134046, 32'sd23611, 32'sd11530, 32'sd954899,
32'sd159524, 32'sd383870, 32'sd73688, 32'sd143562, 32'sd64366, 32'sd946827, 32'sd11797, 32'sd174527, 32'sd275584, 32'sd197917,
32'sd16536, 32'sd34653, 32'sd16574, 32'sd10818, 32'sd207371, 32'sd41463, 32'sd112136, 32'sd358088, 32'sd184645, 32'sd183540,
32'sd558953, 32'sd47295, 32'sd53809, 32'sd77375, 32'sd351827, 32'sd406402, 32'sd345978, 32'sd214617, 32'sd175794, 32'sd152688,
32'sd230075, 32'sd487770, 32'sd283688, 32'sd316757, 32'sd103110, 32'sd144600, 32'sd654875, 32'sd277621, 32'sd390210, 32'sd19230,
32'sd312469, 32'sd93468, 32'sd430210, 32'sd41743, 32'sd206773, 32'sd451031, 32'sd556002, 32'sd595862, 32'sd112300, 32'sd170265,
32'sd164056, 32'sd166572, 32'sd83212, 32'sd477232, 32'sd83002, 32'sd147737, 32'sd366750, 32'sd272816, 32'sd131004, 32'sd234260,
32'sd56574, 32'sd72307, 32'sd109243, 32'sd24332, 32'sd883702, 32'sd308514, 32'sd342533, 32'sd37628, 32'sd32981, 32'sd14829,
32'sd20727, 32'sd27601, 32'sd2236, 32'sd505708, 32'sd367, 32'sd194603, 32'sd560635, 32'sd47421, 32'sd20443, 32'sd495174,
32'sd835489, 32'sd11848, 32'sd89217, 32'sd151949, 32'sd766012, 32'sd7968, 32'sd115197, 32'sd112924, 32'sd590086, 32'sd753100,
32'sd117511, 32'sd396311, 32'sd154850, 32'sd125155, 32'sd80944, 32'sd278981, 32'sd309261, 32'sd145154, 32'sd272387, 32'sd73079,
32'sd262795, 32'sd158210, 32'sd558442, 32'sd42547, 32'sd551056, 32'sd64908, 32'sd10828, 32'sd169245, 32'sd193709, 32'sd20500,
32'sd206937, 32'sd318681, 32'sd752238, 32'sd93711, 32'sd317649, 32'sd23200, 32'sd320962, 32'sd413068, 32'sd646889, 32'sd12784,
32'sd262180, 32'sd192470, 32'sd453316, 32'sd11561, 32'sd483708, 32'sd38000, 32'sd274223, 32'sd411494, 32'sd688816, 32'sd632003,
32'sd384727, 32'sd75310, 32'sd451097, 32'sd193308, 32'sd2990, 32'sd487064, 32'sd75455, 32'sd194045, 32'sd176694, 32'sd167401,
32'sd28482, 32'sd332871, 32'sd20222, 32'sd378777, 32'sd122938, 32'sd148071, 32'sd230046, 32'sd24656, 32'sd447305, 32'sd108780,
32'sd73826, 32'sd64048, 32'sd455611, 32'sd505363, 32'sd697430, 32'sd106091, 32'sd43005, 32'sd218938, 32'sd109756, 32'sd8698,
32'sd323740, 32'sd595962, 32'sd67447, 32'sd335554, 32'sd83882, 32'sd572513, 32'sd530354, 32'sd382100, 32'sd200000, 32'sd50724,
32'sd605867, 32'sd318270, 32'sd74832, 32'sd15510, 32'sd236359, 32'sd187563, 32'sd107160, 32'sd368492, 32'sd152632, 32'sd22941,
32'sd69531, 32'sd42382, 32'sd150714, 32'sd118727, 32'sd410863, 32'sd90792, 32'sd104844, 32'sd9877, 32'sd144363, 32'sd129774,
32'sd100186, 32'sd115297, 32'sd90783, 32'sd830282, 32'sd571529, 32'sd21427, 32'sd279289, 32'sd81594, 32'sd931910, 32'sd204137,
32'sd163823, 32'sd733929, 32'sd190733, 32'sd286413, 32'sd262713, 32'sd238738, 32'sd1881, 32'sd600134, 32'sd145495, 32'sd248985,
32'sd372597, 32'sd244903, 32'sd834960, 32'sd279424, 32'sd44503, 32'sd458166, 32'sd573639, 32'sd156916, 32'sd137415, 32'sd25444,
32'sd71807, 32'sd67420, 32'sd136849, 32'sd624415, 32'sd106442, 32'sd140725, 32'sd244986, 32'sd468852, 32'sd764965, 32'sd185838,
32'sd176452, 32'sd196611, 32'sd62538, 32'sd455113, 32'sd80790, 32'sd259314, 32'sd74867, 32'sd3956, 32'sd189344, 32'sd677448,
32'sd600125, 32'sd776295, 32'sd906659, 32'sd900882, 32'sd55617, 32'sd180478, 32'sd173400, 32'sd437476, 32'sd438780, 32'sd319285,
32'sd561369, 32'sd58675, 32'sd968463, 32'sd61659, 32'sd634713, 32'sd329565, 32'sd209412, 32'sd644436, 32'sd209370, 32'sd326310,
32'sd23565, 32'sd68509, 32'sd130697, 32'sd132276, 32'sd339163, 32'sd253526, 32'sd7941, 32'sd479911, 32'sd356013, 32'sd201632,
32'sd39663, 32'sd558351, 32'sd220716, 32'sd83926, 32'sd263293, 32'sd476402, 32'sd24543, 32'sd19093, 32'sd13736, 32'sd291919,
32'sd49954, 32'sd172708, 32'sd458634, 32'sd254440, 32'sd152164, 32'sd287584, 32'sd22597, 32'sd160179, 32'sd5958, 32'sd42186,
32'sd238547, 32'sd108361, 32'sd29585, 32'sd75182, 32'sd224288, 32'sd834156, 32'sd375899, 32'sd188402, 32'sd518553, 32'sd607336,
32'sd207842, 32'sd32247, 32'sd699288, 32'sd72574, 32'sd59402, 32'sd157320, 32'sd863583, 32'sd195322, 32'sd270694, 32'sd182263,
32'sd158932, 32'sd143030, 32'sd539224, 32'sd4823, 32'sd291930, 32'sd154321, 32'sd217823, 32'sd209724, 32'sd110457, 32'sd3639,
32'sd47671, 32'sd22434, 32'sd212803, 32'sd851506, 32'sd2890, 32'sd204261, 32'sd449197, 32'sd94068, 32'sd548412, 32'sd53505,
32'sd22155, 32'sd45350, 32'sd315133, 32'sd249411, 32'sd34547, 32'sd127519, 32'sd15815, 32'sd131132, 32'sd753951, 32'sd20631,
32'sd65207, 32'sd77716, 32'sd330643, 32'sd54112, 32'sd1689, 32'sd209577, 32'sd604523, 32'sd15442, 32'sd362834, 32'sd744909,
32'sd500422, 32'sd871498, 32'sd53897, 32'sd61377, 32'sd19792, 32'sd637450, 32'sd129165, 32'sd57601, 32'sd83432, 32'sd242650,
32'sd128449, 32'sd60978, 32'sd49271, 32'sd374818, 32'sd804408, 32'sd72072, 32'sd654786, 32'sd59147, 32'sd417296, 32'sd324,
32'sd310933, 32'sd155590, 32'sd77503, 32'sd492286, 32'sd88140, 32'sd109743, 32'sd132496, 32'sd52652, 32'sd169815, 32'sd523232,
32'sd475070, 32'sd63884, 32'sd45312, 32'sd22258, 32'sd938310, 32'sd265396, 32'sd226803, 32'sd150710, 32'sd369930, 32'sd345764,
32'sd75189, 32'sd338897, 32'sd246924, 32'sd34885, 32'sd72446, 32'sd184966, 32'sd228996, 32'sd236647, 32'sd26725, 32'sd17868,
32'sd367998, 32'sd240339, 32'sd95760, 32'sd28860, 32'sd7572, 32'sd162571, 32'sd189930, 32'sd69189, 32'sd30656, 32'sd131771,
32'sd490211, 32'sd350004, 32'sd79368, 32'sd36195, 32'sd129880, 32'sd714150, 32'sd175874, 32'sd41530, 32'sd196567, 32'sd536992,
32'sd684910, 32'sd246010, 32'sd92695, 32'sd216322, 32'sd936956, 32'sd106026, 32'sd790354, 32'sd62814, 32'sd792666, 32'sd67383,
32'sd6274, 32'sd577497, 32'sd235947, 32'sd94637, 32'sd859185, 32'sd214284, 32'sd256282, 32'sd347642, 32'sd449319, 32'sd535918,
32'sd37284, 32'sd8945, 32'sd340421, 32'sd2815, 32'sd233841, 32'sd592079, 32'sd408947, 32'sd13855, 32'sd30827, 32'sd544981,
32'sd130383, 32'sd230925, 32'sd260953, 32'sd15489, 32'sd70335, 32'sd215302, 32'sd29800, 32'sd711459, 32'sd123900, 32'sd755809,
32'sd27278, 32'sd4109, 32'sd342477, 32'sd384920, 32'sd936192, 32'sd39625, 32'sd145036, 32'sd676865, 32'sd315508, 32'sd17882,
32'sd47650, 32'sd101829, 32'sd147061, 32'sd676946, 32'sd363560, 32'sd362798, 32'sd180539, 32'sd520030, 32'sd12829, 32'sd380853,
32'sd53019, 32'sd628976, 32'sd762725, 32'sd229330, 32'sd305736, 32'sd631239, 32'sd463855, 32'sd413061, 32'sd171023, 32'sd441970,
32'sd242858, 32'sd113881, 32'sd64648, 32'sd553112, 32'sd278674, 32'sd69820, 32'sd62415, 32'sd107959, 32'sd458359, 32'sd268421,
32'sd376421, 32'sd311745, 32'sd663631, 32'sd726720, 32'sd394464, 32'sd58156, 32'sd593532, 32'sd148111, 32'sd51429, 32'sd215488,
32'sd186585, 32'sd210465, 32'sd204479, 32'sd200407, 32'sd741033, 32'sd420796, 32'sd260, 32'sd65163, 32'sd1583, 32'sd140244,
32'sd19481, 32'sd308299, 32'sd41578, 32'sd7763, 32'sd182516, 32'sd48012, 32'sd550201, 32'sd34393, 32'sd152360, 32'sd527958,
32'sd147363, 32'sd25696, 32'sd1062706, 32'sd733321, 32'sd22133, 32'sd499056, 32'sd445110, 32'sd364188, 32'sd37268, 32'sd34010,
32'sd14899, 32'sd806278, 32'sd438168, 32'sd194401, 32'sd514615, 32'sd199485, 32'sd206953, 32'sd596155, 32'sd32739, 32'sd478477,
32'sd389323, 32'sd232986, 32'sd43003, 32'sd50132, 32'sd206690, 32'sd393789, 32'sd84667, 32'sd35984, 32'sd402350, 32'sd510442,
32'sd407167, 32'sd637200, 32'sd351812, 32'sd277416, 32'sd171390, 32'sd156876, 32'sd246599, 32'sd304924, 32'sd56427, 32'sd594727,
32'sd28377, 32'sd192383, 32'sd283536, 32'sd93463, 32'sd266448, 32'sd104803, 32'sd29272, 32'sd140594, 32'sd170449, 32'sd6026,
32'sd114241, 32'sd50873, 32'sd180054, 32'sd273349, 32'sd70921, 32'sd270465, 32'sd133597, 32'sd168839, 32'sd56478, 32'sd446486,
32'sd248955, 32'sd108498, 32'sd68230, 32'sd652143, 32'sd134946, 32'sd181801, 32'sd20741, 32'sd20556, 32'sd286007, 32'sd537272,
32'sd178170, 32'sd165361, 32'sd699663, 32'sd212611, 32'sd55669, 32'sd127891, 32'sd191017, 32'sd445351, 32'sd11378, 32'sd35212,
32'sd214136, 32'sd17253, 32'sd264586, 32'sd15561, 32'sd51867, 32'sd131832, 32'sd275370, 32'sd30183, 32'sd52552, 32'sd74796,
32'sd227188, 32'sd469366, 32'sd12631, 32'sd543214, 32'sd225386, 32'sd70158, 32'sd406149, 32'sd314358, 32'sd146192, 32'sd221463,
32'sd22078, 32'sd272813, 32'sd471495, 32'sd18820, 32'sd374620, 32'sd49519, 32'sd569427, 32'sd168650, 32'sd80153, 32'sd267810,
32'sd79411, 32'sd296270, 32'sd111080, 32'sd239794, 32'sd551712, 32'sd163938, 32'sd282028, 32'sd390436, 32'sd386292, 32'sd160444,
32'sd254157, 32'sd46039, 32'sd335337, 32'sd473483, 32'sd169191, 32'sd278230, 32'sd149798, 32'sd11682, 32'sd110581, 32'sd218184,
32'sd141216, 32'sd728850, 32'sd11492, 32'sd460137, 32'sd65553, 32'sd535220, 32'sd626359, 32'sd12878, 32'sd60418, 32'sd435339,
32'sd936045, 32'sd327635, 32'sd781786, 32'sd419798, 32'sd209750, 32'sd148173, 32'sd189941, 32'sd92842, 32'sd141941, 32'sd47700,
32'sd527067, 32'sd123214, 32'sd19078, 32'sd2314, 32'sd626279, 32'sd587203, 32'sd675351, 32'sd209515, 32'sd214165, 32'sd125133,
32'sd82149, 32'sd274731, 32'sd214400, 32'sd54104, 32'sd440053, 32'sd160369, 32'sd99102, 32'sd273594, 32'sd234576, 32'sd208309,
32'sd112322, 32'sd108689, 32'sd354963, 32'sd208823, 32'sd263282, 32'sd41335, 32'sd68117, 32'sd28673, 32'sd365862, 32'sd30550,
32'sd361447, 32'sd241100, 32'sd554997, 32'sd307839, 32'sd331864, 32'sd30311, 32'sd58742, 32'sd413139, 32'sd924733, 32'sd352,
32'sd301785, 32'sd1245402, 32'sd301661, 32'sd116527, 32'sd184800, 32'sd219024, 32'sd106353, 32'sd559919, 32'sd254865, 32'sd50356,
32'sd349077, 32'sd121892, 32'sd27541, 32'sd7248, 32'sd41710, 32'sd50639, 32'sd177017, 32'sd389890, 32'sd322855, 32'sd159681,
32'sd221996, 32'sd296042, 32'sd410103, 32'sd338210, 32'sd411648, 32'sd78529, 32'sd14275, 32'sd62878, 32'sd31295, 32'sd997862,
32'sd22795, 32'sd245133, 32'sd1011088, 32'sd3169, 32'sd407871, 32'sd383211, 32'sd484073, 32'sd276172, 32'sd91488, 32'sd978962,
32'sd183298, 32'sd63346, 32'sd91835, 32'sd521815, 32'sd113068, 32'sd418471, 32'sd35308, 32'sd208478, 32'sd284382, 32'sd795632,
32'sd537591, 32'sd225353, 32'sd404420, 32'sd255744, 32'sd9759, 32'sd196446, 32'sd224603, 32'sd392291, 32'sd241486, 32'sd211397,
32'sd88200, 32'sd659029, 32'sd379550, 32'sd624712, 32'sd602500, 32'sd252379, 32'sd269843, 32'sd56292, 32'sd39505, 32'sd139731,
32'sd71343, 32'sd135662, 32'sd284974, 32'sd393384, 32'sd623131, 32'sd147595, 32'sd43700, 32'sd388254, 32'sd69878, 32'sd54246,
32'sd3215, 32'sd46237, 32'sd26207, 32'sd28803, 32'sd49879, 32'sd49750, 32'sd656677, 32'sd371804, 32'sd180678, 32'sd233551,
32'sd585809, 32'sd391977, 32'sd270810, 32'sd129669, 32'sd922420, 32'sd484252, 32'sd13837, 32'sd75915, 32'sd357097, 32'sd87392,
32'sd348602, 32'sd129501, 32'sd132236, 32'sd1016157, 32'sd58971, 32'sd868873, 32'sd13752, 32'sd217066, 32'sd170576, 32'sd415817,
32'sd597107, 32'sd400174, 32'sd231869, 32'sd618822, 32'sd163362, 32'sd25081, 32'sd152804, 32'sd696021, 32'sd488538, 32'sd1074840,
32'sd249623, 32'sd30440, 32'sd76037, 32'sd365814, 32'sd271038, 32'sd173301, 32'sd458297, 32'sd168449, 32'sd180114, 32'sd33624,
32'sd20667, 32'sd347411, 32'sd715044, 32'sd485753, 32'sd440832, 32'sd164677, 32'sd464024, 32'sd107847, 32'sd250409, 32'sd61896,
32'sd543975, 32'sd62200, 32'sd197098, 32'sd238725, 32'sd805548, 32'sd720970, 32'sd267897, 32'sd708452, 32'sd202151, 32'sd115057,
32'sd344850, 32'sd334525, 32'sd282348, 32'sd620718, 32'sd65388, 32'sd92926, 32'sd675078, 32'sd88350, 32'sd230696, 32'sd238790,
32'sd759559, 32'sd164081, 32'sd80644, 32'sd809336, 32'sd30521, 32'sd103630, 32'sd141455, 32'sd684004, 32'sd317930, 32'sd636191,
32'sd312253, 32'sd198631, 32'sd660085, 32'sd213073, 32'sd476140, 32'sd436666, 32'sd154216, 32'sd871058, 32'sd94219, 32'sd277642,
32'sd95584, 32'sd512396, 32'sd273183, 32'sd691587, 32'sd193478, 32'sd46507, 32'sd286477, 32'sd101741, 32'sd702824, 32'sd222118,
32'sd297004, 32'sd1057720, 32'sd418342, 32'sd548097, 32'sd48768, 32'sd415108, 32'sd18292, 32'sd8525, 32'sd38362, 32'sd344237,
32'sd213639, 32'sd58119, 32'sd65593, 32'sd200458, 32'sd375187, 32'sd136439, 32'sd214763, 32'sd47022, 32'sd122682, 32'sd61134,
32'sd19460, 32'sd59091, 32'sd144046, 32'sd357474, 32'sd566513, 32'sd671137, 32'sd326541, 32'sd529528, 32'sd660163, 32'sd147721,
32'sd122351, 32'sd541554, 32'sd247956, 32'sd282780, 32'sd488228, 32'sd285346, 32'sd77916, 32'sd74456, 32'sd11256, 32'sd494934,
32'sd238920, 32'sd483111, 32'sd269979, 32'sd9742, 32'sd656412, 32'sd92154, 32'sd213984, 32'sd1076930, 32'sd29863, 32'sd366757,
32'sd148543, 32'sd115211, 32'sd551956, 32'sd107439, 32'sd444607, 32'sd73510, 32'sd58460, 32'sd66778, 32'sd284199, 32'sd172706,
32'sd104431, 32'sd50350, 32'sd359739, 32'sd107392, 32'sd76423, 32'sd181620, 32'sd416883, 32'sd877577, 32'sd342380, 32'sd645785,
32'sd131993, 32'sd711508, 32'sd85683, 32'sd36457, 32'sd77866, 32'sd67251, 32'sd441510, 32'sd20564, 32'sd180406, 32'sd834385,
32'sd96879, 32'sd435362, 32'sd39232, 32'sd111171, 32'sd273924, 32'sd29474, 32'sd786640, 32'sd16908, 32'sd601518, 32'sd10620,
32'sd5273, 32'sd194599, 32'sd366019, 32'sd35657, 32'sd535437, 32'sd514007, 32'sd8491, 32'sd753858, 32'sd100337, 32'sd213685,
32'sd21870, 32'sd514143, 32'sd23355, 32'sd468270, 32'sd72524, 32'sd726338, 32'sd292207, 32'sd72250, 32'sd323669, 32'sd539506,
32'sd9899, 32'sd70052, 32'sd657182, 32'sd92451, 32'sd156067, 32'sd54816, 32'sd164187, 32'sd246168, 32'sd294910, 32'sd142897,
32'sd227643, 32'sd29767, 32'sd381073, 32'sd136387, 32'sd105426, 32'sd549131, 32'sd236567, 32'sd98461, 32'sd94284, 32'sd9774,
32'sd12827, 32'sd43381, 32'sd355813, 32'sd191698, 32'sd114838, 32'sd34095, 32'sd127904, 32'sd595579, 32'sd12683, 32'sd490889,
32'sd42211, 32'sd743028, 32'sd23219, 32'sd483321, 32'sd473901, 32'sd236242, 32'sd252968, 32'sd434715, 32'sd72813, 32'sd200025,
32'sd241002, 32'sd184919, 32'sd146174, 32'sd79921, 32'sd55308, 32'sd520058, 32'sd263799, 32'sd268597, 32'sd219050, 32'sd177846,
32'sd418811, 32'sd434203, 32'sd311436, 32'sd167826, 32'sd175468, 32'sd321126, 32'sd177949, 32'sd90591, 32'sd468802, 32'sd652339,
32'sd529204, 32'sd412678, 32'sd132010, 32'sd126409, 32'sd414356, 32'sd371934, 32'sd296097, 32'sd83105, 32'sd192659, 32'sd173456,
32'sd113325, 32'sd100289, 32'sd364874, 32'sd232363, 32'sd34469, 32'sd428501, 32'sd274826, 32'sd67299, 32'sd3727, 32'sd965498,
32'sd117957, 32'sd346425, 32'sd110988, 32'sd43780, 32'sd616086, 32'sd1173499, 32'sd66284, 32'sd54513, 32'sd98943, 32'sd382633,
32'sd233222, 32'sd39193, 32'sd48160, 32'sd232203, 32'sd146285, 32'sd635555, 32'sd120734, 32'sd2067, 32'sd22612, 32'sd159415,
32'sd123548, 32'sd188140, 32'sd318894, 32'sd117745, 32'sd52712, 32'sd65562, 32'sd48211, 32'sd215360, 32'sd643934, 32'sd127675,
32'sd544766, 32'sd190788, 32'sd143615, 32'sd584037, 32'sd390683, 32'sd193172, 32'sd792930, 32'sd408093, 32'sd283783, 32'sd4878,
32'sd12580, 32'sd304183, 32'sd82042, 32'sd97822, 32'sd661815, 32'sd44941, 32'sd742888, 32'sd325692, 32'sd287678, 32'sd416110,
32'sd171673, 32'sd280794, 32'sd289426, 32'sd45847, 32'sd116599, 32'sd425488, 32'sd199263, 32'sd117846, 32'sd170933, 32'sd282061,
32'sd633180, 32'sd160478, 32'sd69303, 32'sd1158637, 32'sd22008, 32'sd155918, 32'sd643282, 32'sd316115, 32'sd361252, 32'sd168862,
32'sd319548, 32'sd330089, 32'sd422759, 32'sd178848, 32'sd160995, 32'sd730569, 32'sd320492, 32'sd435823, 32'sd98161, 32'sd109799,
32'sd106705, 32'sd153513, 32'sd182247, 32'sd405889, 32'sd90468, 32'sd164081, 32'sd330080, 32'sd201669, 32'sd128716, 32'sd420048,
32'sd33820, 32'sd188758, 32'sd857776, 32'sd298595, 32'sd187455, 32'sd234151, 32'sd376351, 32'sd460685, 32'sd716068, 32'sd278741,
32'sd139774, 32'sd366667, 32'sd130474, 32'sd319458, 32'sd116963, 32'sd266009, 32'sd235051, 32'sd170341, 32'sd557043, 32'sd185347,
32'sd137854, 32'sd9493, 32'sd383939, 32'sd100177, 32'sd7041, 32'sd129794, 32'sd52063, 32'sd755020, 32'sd1019235, 32'sd428462,
32'sd549703, 32'sd244245, 32'sd16565, 32'sd79193, 32'sd937453, 32'sd1343153, 32'sd47443, 32'sd1078090, 32'sd161980, 32'sd336013,
32'sd479084, 32'sd377949, 32'sd164277, 32'sd128234, 32'sd170328, 32'sd108723, 32'sd8218, 32'sd119884, 32'sd150997, 32'sd96841,
32'sd180748, 32'sd99360, 32'sd719124, 32'sd302399, 32'sd787, 32'sd427089, 32'sd359782, 32'sd70944, 32'sd97659, 32'sd21997,
32'sd65476, 32'sd50515, 32'sd968391, 32'sd21881, 32'sd118754, 32'sd486271, 32'sd30768, 32'sd32504, 32'sd359509, 32'sd698394,
32'sd208837, 32'sd265149, 32'sd83576, 32'sd92461, 32'sd5891, 32'sd338198, 32'sd418603, 32'sd18112, 32'sd435237, 32'sd60434,
32'sd95626, 32'sd567330, 32'sd24458, 32'sd350641, 32'sd21778, 32'sd74850, 32'sd80522, 32'sd90195, 32'sd119824, 32'sd342993,
32'sd93751, 32'sd187236, 32'sd30065, 32'sd448662, 32'sd91949, 32'sd321224, 32'sd16433, 32'sd38347, 32'sd20473, 32'sd221882,
32'sd3986, 32'sd461875, 32'sd536551, 32'sd4446, 32'sd839678, 32'sd509716, 32'sd26214, 32'sd677242, 32'sd121000, 32'sd192780,
32'sd905601, 32'sd305329, 32'sd56745, 32'sd473561, 32'sd506760, 32'sd388720, 32'sd16146, 32'sd325458, 32'sd705170, 32'sd26366,
32'sd237319, 32'sd136543, 32'sd98124, 32'sd316090, 32'sd17513, 32'sd250928, 32'sd48798, 32'sd129622, 32'sd136605, 32'sd231514,
32'sd240356, 32'sd110036, 32'sd546168, 32'sd151711, 32'sd165860, 32'sd345381, 32'sd36714, 32'sd280016, 32'sd132272, 32'sd97546,
32'sd338572, 32'sd17095, 32'sd434541, 32'sd111911, 32'sd387076, 32'sd592391, 32'sd443034, 32'sd430138, 32'sd102716, 32'sd612953,
32'sd97844, 32'sd210416, 32'sd490859, 32'sd108195, 32'sd101849, 32'sd813753, 32'sd317752, 32'sd168992, 32'sd438861, 32'sd158866,
32'sd632151, 32'sd235353, 32'sd101874, 32'sd244518, 32'sd541395, 32'sd787072, 32'sd352677, 32'sd452299, 32'sd29305, 32'sd254726,
32'sd13173, 32'sd598046, 32'sd42386, 32'sd731764, 32'sd186090, 32'sd152620, 32'sd694190, 32'sd154552, 32'sd13935, 32'sd249679,
32'sd374185, 32'sd92125, 32'sd71121, 32'sd43641, 32'sd587536, 32'sd242297, 32'sd30745, 32'sd91902, 32'sd131842, 32'sd638675,
32'sd77317, 32'sd692025, 32'sd121666, 32'sd483951, 32'sd23456, 32'sd227821, 32'sd582545, 32'sd39204, 32'sd285268, 32'sd1036525,
32'sd206948, 32'sd206500, 32'sd31290, 32'sd529890, 32'sd104705, 32'sd246046, 32'sd340640, 32'sd656953, 32'sd378520, 32'sd115183,
32'sd362202, 32'sd199431, 32'sd175695, 32'sd291750, 32'sd141980, 32'sd14713, 32'sd196479, 32'sd31121, 32'sd221602, 32'sd958083,
32'sd350782, 32'sd454277, 32'sd721505, 32'sd391210, 32'sd1800, 32'sd45304, 32'sd131103, 32'sd171536, 32'sd309956, 32'sd1200013,
32'sd186492, 32'sd73925, 32'sd66162, 32'sd61088, 32'sd128951, 32'sd5032, 32'sd313072, 32'sd128839, 32'sd6284, 32'sd78303,
32'sd602268, 32'sd50043, 32'sd1451115, 32'sd477797, 32'sd20852, 32'sd175084, 32'sd166808, 32'sd345917, 32'sd352657, 32'sd566587,
32'sd268985, 32'sd7181, 32'sd472398, 32'sd144388, 32'sd212321, 32'sd841247, 32'sd28415, 32'sd5976, 32'sd49362, 32'sd436290,
32'sd582499, 32'sd1028190, 32'sd293666, 32'sd224386, 32'sd94557, 32'sd160636, 32'sd593307, 32'sd228204, 32'sd48298, 32'sd350883,
32'sd45916, 32'sd262199, 32'sd316127, 32'sd91756, 32'sd116174, 32'sd269293, 32'sd362972, 32'sd156894, 32'sd666004, 32'sd218395,
32'sd13363, 32'sd22934, 32'sd244228, 32'sd66065, 32'sd121941, 32'sd147152, 32'sd503872, 32'sd675752, 32'sd269407, 32'sd209139,
32'sd95856, 32'sd5826, 32'sd13213, 32'sd405074, 32'sd276331, 32'sd164677, 32'sd57315, 32'sd113152, 32'sd72636, 32'sd121623,
32'sd43236, 32'sd426151, 32'sd154316, 32'sd183897, 32'sd258850, 32'sd27486, 32'sd51308, 32'sd98190, 32'sd130994, 32'sd77207,
32'sd327046, 32'sd512037, 32'sd272165, 32'sd380690, 32'sd214280, 32'sd835420, 32'sd406880, 32'sd63444, 32'sd675235, 32'sd419097,
32'sd585352, 32'sd440227, 32'sd259936, 32'sd693634, 32'sd468214, 32'sd298364, 32'sd118316, 32'sd227218, 32'sd217684, 32'sd273397,
32'sd105906, 32'sd557700, 32'sd28048, 32'sd399004, 32'sd207778, 32'sd56878, 32'sd288370, 32'sd216027, 32'sd483574, 32'sd375676,
32'sd280320, 32'sd532973, 32'sd24802, 32'sd27727, 32'sd50356, 32'sd524622, 32'sd277122, 32'sd188435, 32'sd109250, 32'sd773598,
32'sd452827, 32'sd193599, 32'sd185268, 32'sd404339, 32'sd89071, 32'sd276666, 32'sd277348, 32'sd188710, 32'sd863431, 32'sd409437,
32'sd238909, 32'sd225364, 32'sd345707, 32'sd161982, 32'sd242907, 32'sd204, 32'sd1292290, 32'sd183043, 32'sd39382, 32'sd32675,
32'sd233367, 32'sd164049, 32'sd1048553, 32'sd130651, 32'sd956698, 32'sd86006, 32'sd162039, 32'sd223030, 32'sd184320, 32'sd67705,
32'sd6618, 32'sd118161, 32'sd138760, 32'sd1064989, 32'sd118308, 32'sd223165, 32'sd491931, 32'sd100344, 32'sd18033, 32'sd66583,
32'sd188137, 32'sd309120, 32'sd556707, 32'sd103689, 32'sd244351, 32'sd60718, 32'sd613056, 32'sd54321, 32'sd359841, 32'sd38486,
32'sd298612, 32'sd706156, 32'sd84096, 32'sd226016, 32'sd29527, 32'sd54589, 32'sd29975, 32'sd1109504, 32'sd137232, 32'sd880103,
32'sd64896, 32'sd553485, 32'sd170813, 32'sd34358, 32'sd82974, 32'sd324731, 32'sd73514, 32'sd458216, 32'sd203058, 32'sd2670,
32'sd125880, 32'sd305354, 32'sd729793, 32'sd54977, 32'sd177586, 32'sd479798, 32'sd303228, 32'sd440380, 32'sd147199, 32'sd348333,
32'sd170373, 32'sd251696, 32'sd163550, 32'sd578520, 32'sd1232687, 32'sd25780, 32'sd347423, 32'sd379568, 32'sd506744, 32'sd117027,
32'sd410990, 32'sd50523, 32'sd30273, 32'sd98248, 32'sd129387, 32'sd89639, 32'sd690001, 32'sd103029, 32'sd108862, 32'sd165928,
32'sd872343, 32'sd1269723, 32'sd40395, 32'sd191952, 32'sd351661, 32'sd560568, 32'sd287719, 32'sd292268, 32'sd349465, 32'sd238894,
32'sd17649, 32'sd358529, 32'sd303720, 32'sd351697, 32'sd22416, 32'sd564940, 32'sd283204, 32'sd361786, 32'sd181648, 32'sd367204,
32'sd61194, 32'sd263279, 32'sd182598, 32'sd208154, 32'sd82452, 32'sd684121, 32'sd248647, 32'sd9625, 32'sd69489, 32'sd444977,
32'sd625984, 32'sd176027, 32'sd171632, 32'sd329243, 32'sd40557, 32'sd482206, 32'sd571774, 32'sd289030, 32'sd30643, 32'sd676227,
32'sd532018, 32'sd86844, 32'sd120692, 32'sd125443, 32'sd209255, 32'sd443988, 32'sd148920, 32'sd1190841, 32'sd1044122, 32'sd131149,
32'sd70916, 32'sd16088, 32'sd312464, 32'sd241109, 32'sd866339, 32'sd33852, 32'sd14677, 32'sd142965, 32'sd56572, 32'sd78720,
32'sd79323, 32'sd148599, 32'sd169816, 32'sd126783, 32'sd363354, 32'sd95143, 32'sd6716, 32'sd326386, 32'sd323649, 32'sd393392,
32'sd310455, 32'sd181260, 32'sd340461, 32'sd626962, 32'sd728082, 32'sd600495, 32'sd337058, 32'sd93171, 32'sd72579, 32'sd309076,
32'sd180182, 32'sd466241, 32'sd446744, 32'sd33106, 32'sd289864, 32'sd57647, 32'sd392952, 32'sd509257, 32'sd89292, 32'sd153508,
32'sd236351, 32'sd38285, 32'sd82495, 32'sd688411, 32'sd649964, 32'sd438215, 32'sd205597, 32'sd549589, 32'sd391209, 32'sd473595,
32'sd780551, 32'sd178934, 32'sd781665, 32'sd348252, 32'sd25825, 32'sd105698, 32'sd124532, 32'sd110039, 32'sd154504, 32'sd521170,
32'sd10530, 32'sd707334, 32'sd755833, 32'sd453158, 32'sd344287, 32'sd297791, 32'sd111472, 32'sd234386, 32'sd67386, 32'sd578704,
32'sd14783, 32'sd139181, 32'sd497884, 32'sd60377, 32'sd5644, 32'sd123532, 32'sd38645, 32'sd538991, 32'sd275597, 32'sd210496,
32'sd246960, 32'sd46062, 32'sd68889, 32'sd545460, 32'sd203593, 32'sd519307, 32'sd86514, 32'sd170152, 32'sd6190, 32'sd10109,
32'sd408544, 32'sd247881, 32'sd159694, 32'sd42081, 32'sd148333, 32'sd234156, 32'sd67504, 32'sd131148, 32'sd167612, 32'sd18991,
32'sd387696, 32'sd85415, 32'sd479362, 32'sd146740, 32'sd3242, 32'sd278563, 32'sd61537, 32'sd135324, 32'sd31773, 32'sd78547,
32'sd638003, 32'sd327757, 32'sd65594, 32'sd387827, 32'sd230626, 32'sd370689, 32'sd246803, 32'sd137475, 32'sd41062, 32'sd370355,
32'sd29082, 32'sd324553, 32'sd59418, 32'sd542516, 32'sd879275, 32'sd379285, 32'sd689703, 32'sd250040, 32'sd5708, 32'sd576175,
32'sd208187, 32'sd186298, 32'sd895491, 32'sd790109, 32'sd149130, 32'sd300792, 32'sd559411, 32'sd729703, 32'sd869530, 32'sd965487,
32'sd237789, 32'sd241520, 32'sd604519, 32'sd112724, 32'sd1406, 32'sd344028, 32'sd410826, 32'sd44841, 32'sd401933, 32'sd599203,
32'sd54231, 32'sd13261, 32'sd219132, 32'sd54657, 32'sd24312, 32'sd189901, 32'sd364050, 32'sd88878, 32'sd194033, 32'sd493108,
32'sd608752, 32'sd226918, 32'sd15262, 32'sd515662, 32'sd257721, 32'sd267162, 32'sd52432, 32'sd321629, 32'sd8767, 32'sd418285,
32'sd47880, 32'sd517052, 32'sd22494, 32'sd857530, 32'sd103367, 32'sd203538, 32'sd151544, 32'sd532659, 32'sd615524, 32'sd220892,
32'sd310779, 32'sd173591, 32'sd48852, 32'sd266098, 32'sd40935, 32'sd23125, 32'sd28386, 32'sd99543, 32'sd75792, 32'sd287896,
32'sd149488, 32'sd250373, 32'sd162992, 32'sd88057, 32'sd38919, 32'sd528112, 32'sd373441, 32'sd596905, 32'sd555478, 32'sd18880,
32'sd232530, 32'sd23029, 32'sd268801, 32'sd331642, 32'sd221538, 32'sd136800, 32'sd145200, 32'sd444488, 32'sd9747, 32'sd105019,
32'sd233993, 32'sd155629, 32'sd225225, 32'sd218301, 32'sd48782, 32'sd196476, 32'sd323892, 32'sd301831, 32'sd497968, 32'sd443383,
32'sd94043, 32'sd769155, 32'sd35286, 32'sd508981, 32'sd69748, 32'sd533385, 32'sd21781, 32'sd191328, 32'sd211020, 32'sd185031,
32'sd794737, 32'sd61042, 32'sd407204, 32'sd636729, 32'sd70125, 32'sd396520, 32'sd688494, 32'sd170231, 32'sd181887, 32'sd239949,
32'sd69457, 32'sd554501, 32'sd312939, 32'sd320629, 32'sd391843, 32'sd280338, 32'sd78602, 32'sd355279, 32'sd1148561, 32'sd128763,
32'sd546079, 32'sd18448, 32'sd166105, 32'sd632269, 32'sd302578, 32'sd1242669, 32'sd947106, 32'sd569746, 32'sd295451, 32'sd66552,
32'sd972264, 32'sd189872, 32'sd3877, 32'sd169238, 32'sd54782, 32'sd84015, 32'sd234780, 32'sd116708, 32'sd351709, 32'sd274417,
32'sd179394, 32'sd344362, 32'sd592293, 32'sd318380, 32'sd54456, 32'sd67537, 32'sd215557, 32'sd102746, 32'sd108639, 32'sd564670,
32'sd76221, 32'sd264517, 32'sd465510, 32'sd119209, 32'sd244435, 32'sd121088, 32'sd261758, 32'sd761100, 32'sd84352, 32'sd626929,
32'sd24979, 32'sd111719, 32'sd371115, 32'sd148398, 32'sd699664, 32'sd429729, 32'sd10086, 32'sd79085, 32'sd734, 32'sd892938,
32'sd108338, 32'sd397110, 32'sd406367, 32'sd234562, 32'sd140251, 32'sd517712, 32'sd69712, 32'sd36615, 32'sd7829, 32'sd626125,
32'sd190920, 32'sd52999, 32'sd989678, 32'sd165369, 32'sd186816, 32'sd605305, 32'sd612452, 32'sd580216, 32'sd99817, 32'sd2297,
32'sd1386506, 32'sd17246, 32'sd111462, 32'sd395525, 32'sd406823, 32'sd91967, 32'sd48731, 32'sd114275, 32'sd1602, 32'sd15225,
32'sd138863, 32'sd82013, 32'sd587371, 32'sd317071, 32'sd42041, 32'sd54524, 32'sd115684, 32'sd65372, 32'sd115587, 32'sd101912,
32'sd177599, 32'sd324, 32'sd147085, 32'sd151377, 32'sd341654, 32'sd490260, 32'sd167156, 32'sd482889, 32'sd351639, 32'sd73723,
32'sd144431, 32'sd87916, 32'sd139365, 32'sd90437, 32'sd137915, 32'sd441056, 32'sd137376, 32'sd346624, 32'sd362740, 32'sd300701,
32'sd199205, 32'sd316883, 32'sd1065515, 32'sd221770, 32'sd205184, 32'sd7801, 32'sd175887, 32'sd94366, 32'sd111332, 32'sd36113,
32'sd364904, 32'sd34238, 32'sd313789, 32'sd206972, 32'sd255027, 32'sd681447, 32'sd123959, 32'sd363328, 32'sd454596, 32'sd23100,
32'sd345301, 32'sd117819, 32'sd878454, 32'sd98411, 32'sd404899, 32'sd203986, 32'sd359271, 32'sd180797, 32'sd156774, 32'sd99873,
32'sd437118, 32'sd112356, 32'sd128804, 32'sd422832, 32'sd694025, 32'sd157732, 32'sd76544, 32'sd145308, 32'sd278053, 32'sd659970,
32'sd49317, 32'sd76246, 32'sd701486, 32'sd752880, 32'sd538317, 32'sd22373, 32'sd86532, 32'sd169758, 32'sd520822, 32'sd2895,
32'sd238623, 32'sd528372, 32'sd232206, 32'sd479843, 32'sd52668, 32'sd66728, 32'sd293748, 32'sd535324, 32'sd230634, 32'sd21496,
32'sd318229, 32'sd267340, 32'sd209747, 32'sd28974, 32'sd252078, 32'sd670482, 32'sd1176795, 32'sd430819, 32'sd438317, 32'sd160237,
32'sd1086, 32'sd192516, 32'sd1270732, 32'sd1109244, 32'sd122434, 32'sd1075655, 32'sd99374, 32'sd388918, 32'sd91219, 32'sd467195,
32'sd51322, 32'sd218585, 32'sd320612, 32'sd29664, 32'sd34852, 32'sd546102, 32'sd36322, 32'sd324696, 32'sd283540, 32'sd2987,
32'sd323419, 32'sd47385, 32'sd428402, 32'sd637491, 32'sd99588, 32'sd482415, 32'sd53177, 32'sd39964, 32'sd542016, 32'sd639242,
32'sd502402, 32'sd1272499, 32'sd123510, 32'sd210281, 32'sd605458, 32'sd629600, 32'sd73471, 32'sd500657, 32'sd354955, 32'sd18271,
32'sd192056, 32'sd21403, 32'sd207104, 32'sd64321, 32'sd46288, 32'sd7920, 32'sd471199, 32'sd14308, 32'sd25119, 32'sd37514,
32'sd61130, 32'sd264025, 32'sd829833, 32'sd225676, 32'sd176240, 32'sd104568, 32'sd517875, 32'sd54529, 32'sd955670, 32'sd70056,
32'sd184510, 32'sd62265, 32'sd513115, 32'sd232154, 32'sd680363, 32'sd561986, 32'sd451891, 32'sd1505510, 32'sd564259, 32'sd54640,
32'sd3821, 32'sd145588, 32'sd44827, 32'sd406228, 32'sd329923, 32'sd255818, 32'sd53867, 32'sd882367, 32'sd786092, 32'sd704081,
32'sd133290, 32'sd346962, 32'sd627265, 32'sd784160, 32'sd211615, 32'sd720007, 32'sd137294, 32'sd101686, 32'sd59026, 32'sd115400,
32'sd528660, 32'sd1017382, 32'sd10488, 32'sd71451, 32'sd11325, 32'sd121254, 32'sd152875, 32'sd30298, 32'sd74742, 32'sd91962,
32'sd701859, 32'sd435259, 32'sd140557, 32'sd199599, 32'sd35550, 32'sd24045, 32'sd647743, 32'sd65698, 32'sd1064920, 32'sd827416,
32'sd308685, 32'sd122223, 32'sd323141, 32'sd244352, 32'sd359440, 32'sd380238, 32'sd16870, 32'sd333872, 32'sd245696, 32'sd261400,
32'sd274779, 32'sd44844, 32'sd265221, 32'sd396078, 32'sd80620, 32'sd184478, 32'sd667074, 32'sd980979, 32'sd401426, 32'sd200626,
32'sd112464, 32'sd518, 32'sd922231, 32'sd392052, 32'sd311908, 32'sd93686, 32'sd157480, 32'sd354537, 32'sd251911, 32'sd176722,
32'sd219720, 32'sd216347, 32'sd157198, 32'sd48950, 32'sd511610, 32'sd160415, 32'sd15595, 32'sd1246374, 32'sd476153, 32'sd65196,
32'sd164217, 32'sd282850, 32'sd726154, 32'sd313437, 32'sd363849, 32'sd113740, 32'sd96219, 32'sd575473, 32'sd28826, 32'sd316771,
32'sd327733, 32'sd34398, 32'sd209446, 32'sd29828, 32'sd444891, 32'sd92618, 32'sd232726, 32'sd734842, 32'sd653069, 32'sd6310,
32'sd937419, 32'sd63, 32'sd181623, 32'sd33509, 32'sd4910, 32'sd53657, 32'sd101372, 32'sd82272, 32'sd82368, 32'sd256083,
32'sd445505, 32'sd167389, 32'sd202897, 32'sd165618, 32'sd650692, 32'sd643203, 32'sd182217, 32'sd338513, 32'sd318163, 32'sd664243,
32'sd406004, 32'sd7084, 32'sd319200, 32'sd192102, 32'sd971908, 32'sd655159, 32'sd667790, 32'sd702202, 32'sd136126, 32'sd197760,
32'sd423185, 32'sd24303, 32'sd63261, 32'sd168754, 32'sd75008, 32'sd4080, 32'sd52405, 32'sd47445, 32'sd41976, 32'sd270280,
32'sd500515, 32'sd14864, 32'sd20237, 32'sd118697, 32'sd216773, 32'sd63456, 32'sd134208, 32'sd444215, 32'sd69548, 32'sd47385,
32'sd1264585, 32'sd46282, 32'sd204762, 32'sd108328, 32'sd47443, 32'sd421143, 32'sd288111, 32'sd469135, 32'sd295436, 32'sd365277,
32'sd28215, 32'sd242463, 32'sd692662, 32'sd83396, 32'sd173153, 32'sd113241, 32'sd7004, 32'sd187731, 32'sd39087, 32'sd239620,
32'sd259981, 32'sd205159, 32'sd226269, 32'sd633, 32'sd446767, 32'sd79362, 32'sd537498, 32'sd148308, 32'sd663019, 32'sd509765,
32'sd196157, 32'sd69352, 32'sd186597, 32'sd367281, 32'sd38623, 32'sd15781, 32'sd95290, 32'sd194036, 32'sd454410, 32'sd50073,
32'sd374602, 32'sd189481, 32'sd123917, 32'sd656242, 32'sd594890, 32'sd157868, 32'sd580365, 32'sd372014, 32'sd111628, 32'sd471797,
32'sd120729, 32'sd837041, 32'sd249644, 32'sd676468, 32'sd161437, 32'sd451169, 32'sd40094, 32'sd634351, 32'sd209746, 32'sd6251,
32'sd91920, 32'sd231178, 32'sd604257, 32'sd974387, 32'sd203434, 32'sd45974, 32'sd4422, 32'sd584284, 32'sd348024, 32'sd9337,
32'sd618846, 32'sd134351, 32'sd461518, 32'sd92884, 32'sd70210, 32'sd382434, 32'sd17649, 32'sd34703, 32'sd243896, 32'sd263250,
32'sd249617, 32'sd228341, 32'sd392629, 32'sd159622, 32'sd416564, 32'sd135192, 32'sd181864, 32'sd553825, 32'sd115593, 32'sd226569,
32'sd641147, 32'sd26854, 32'sd89391, 32'sd64659, 32'sd274419, 32'sd218630, 32'sd895197, 32'sd186205, 32'sd82295, 32'sd388119,
32'sd359510, 32'sd472780, 32'sd319364, 32'sd49544, 32'sd1108930, 32'sd73740, 32'sd63568, 32'sd345561, 32'sd343876, 32'sd17830,
32'sd791, 32'sd197960, 32'sd29516, 32'sd433803, 32'sd9497, 32'sd605412, 32'sd196900, 32'sd436678, 32'sd473055, 32'sd465445,
32'sd147953, 32'sd349683, 32'sd220262, 32'sd476068, 32'sd20982, 32'sd85219, 32'sd423015, 32'sd123336, 32'sd107333, 32'sd34034,
32'sd323204, 32'sd324007, 32'sd367289, 32'sd121344, 32'sd308951, 32'sd111506, 32'sd724467, 32'sd39663, 32'sd367266, 32'sd315525,
32'sd219203, 32'sd55625, 32'sd128953, 32'sd134352, 32'sd688476, 32'sd246597, 32'sd606596, 32'sd387889, 32'sd515484, 32'sd42984,
32'sd439327, 32'sd220623, 32'sd206944, 32'sd188003, 32'sd835069, 32'sd231775, 32'sd54063, 32'sd37760, 32'sd71715, 32'sd212184,
32'sd341444, 32'sd145606, 32'sd15722, 32'sd47658, 32'sd473537, 32'sd192944, 32'sd263336, 32'sd608167, 32'sd90334, 32'sd244524,
32'sd222647, 32'sd346850, 32'sd91785, 32'sd515579, 32'sd750143, 32'sd246270, 32'sd69342, 32'sd491745, 32'sd684666, 32'sd135270,
32'sd472128, 32'sd229534, 32'sd147981, 32'sd87724, 32'sd592358, 32'sd511005, 32'sd65832, 32'sd254791, 32'sd370566, 32'sd471677,
32'sd88014, 32'sd51407, 32'sd162386, 32'sd69300, 32'sd92757, 32'sd191940, 32'sd47115, 32'sd422380, 32'sd88063, 32'sd591215,
32'sd776288, 32'sd311320, 32'sd257620, 32'sd595509, 32'sd209431, 32'sd573070, 32'sd55106, 32'sd227236, 32'sd127288, 32'sd347520,
32'sd186335, 32'sd382248, 32'sd358683, 32'sd70416, 32'sd112155, 32'sd778231, 32'sd237283, 32'sd555572, 32'sd182804, 32'sd415399,
32'sd92600, 32'sd43266, 32'sd680789, 32'sd225339, 32'sd420288, 32'sd474404, 32'sd163838, 32'sd311174, 32'sd703443, 32'sd204763,
32'sd281408, 32'sd447879, 32'sd683323, 32'sd417779, 32'sd229617, 32'sd812651, 32'sd476134, 32'sd87827, 32'sd272930, 32'sd325066,
32'sd247023, 32'sd114766, 32'sd315287, 32'sd301417, 32'sd292876, 32'sd297773, 32'sd152574, 32'sd51717, 32'sd47532, 32'sd227617,
32'sd107188, 32'sd679352, 32'sd70347, 32'sd52902, 32'sd448842, 32'sd619892, 32'sd374031, 32'sd178119, 32'sd222054, 32'sd308904,
32'sd205112, 32'sd60195, 32'sd219248, 32'sd51308, 32'sd211674, 32'sd155466, 32'sd101008, 32'sd218973, 32'sd59755, 32'sd11117,
32'sd393099, 32'sd73437, 32'sd33713, 32'sd434201, 32'sd264930, 32'sd581485, 32'sd5604, 32'sd615499, 32'sd62239, 32'sd104473,
32'sd102898, 32'sd66459, 32'sd154339, 32'sd46954, 32'sd288319, 32'sd671389, 32'sd128205, 32'sd45251, 32'sd137569, 32'sd1130,
32'sd158245, 32'sd39285, 32'sd464176, 32'sd82470, 32'sd660840, 32'sd596090, 32'sd267055, 32'sd143231, 32'sd194929, 32'sd20862,
32'sd588599, 32'sd288696, 32'sd324753, 32'sd76469, 32'sd478072, 32'sd531847, 32'sd86826, 32'sd496258, 32'sd113090, 32'sd525035,
32'sd697090, 32'sd325769, 32'sd76595, 32'sd59129, 32'sd283994, 32'sd113493, 32'sd331398, 32'sd201024, 32'sd566264, 32'sd829642,
32'sd170206, 32'sd91886, 32'sd409205, 32'sd10681, 32'sd553668, 32'sd116935, 32'sd311948, 32'sd944122, 32'sd56010, 32'sd413749,
32'sd153283, 32'sd364248, 32'sd64503, 32'sd239223, 32'sd221545, 32'sd410803, 32'sd57254, 32'sd19971, 32'sd546952, 32'sd36520,
32'sd226268, 32'sd602808, 32'sd116512, 32'sd42909, 32'sd153986, 32'sd178815, 32'sd185577, 32'sd221704, 32'sd278751, 32'sd394001,
32'sd531378, 32'sd50448, 32'sd54609, 32'sd508398, 32'sd28640, 32'sd432100, 32'sd92870, 32'sd103096, 32'sd23623, 32'sd240487,
32'sd192641, 32'sd552493, 32'sd111155, 32'sd384616, 32'sd1144230, 32'sd206935, 32'sd44227, 32'sd570550, 32'sd78624, 32'sd144739,
32'sd301264, 32'sd189543, 32'sd192993, 32'sd361565, 32'sd614209, 32'sd858964, 32'sd233066, 32'sd416857, 32'sd104874, 32'sd521577,
32'sd440960, 32'sd165154, 32'sd16541, 32'sd256337, 32'sd291811, 32'sd8046, 32'sd431009, 32'sd432757, 32'sd381947, 32'sd108161,
32'sd337589, 32'sd288365, 32'sd112648, 32'sd114694, 32'sd82104, 32'sd42074, 32'sd86337, 32'sd346845, 32'sd127584, 32'sd500263,
32'sd140976, 32'sd590871, 32'sd315877, 32'sd24612, 32'sd50321, 32'sd418760, 32'sd38460, 32'sd225986, 32'sd249475, 32'sd68856,
32'sd27706, 32'sd109252, 32'sd348998, 32'sd156842, 32'sd636582, 32'sd48111, 32'sd828396, 32'sd75666, 32'sd63794, 32'sd217800,
32'sd449271, 32'sd188549, 32'sd22067, 32'sd248777, 32'sd490656, 32'sd138377, 32'sd244620, 32'sd73484, 32'sd153933, 32'sd366651,
32'sd30289, 32'sd634991, 32'sd4935, 32'sd971036, 32'sd93837, 32'sd650419, 32'sd152958, 32'sd107450, 32'sd21092, 32'sd960672,
32'sd424872, 32'sd178694, 32'sd7396, 32'sd112100, 32'sd280474, 32'sd68971, 32'sd167466, 32'sd654514, 32'sd253830, 32'sd158990,
32'sd99276, 32'sd3586, 32'sd69354, 32'sd872019, 32'sd639116, 32'sd79660, 32'sd36566, 32'sd247034, 32'sd684971, 32'sd248973,
32'sd291961, 32'sd512157, 32'sd82369, 32'sd692077, 32'sd342622, 32'sd168804, 32'sd44867, 32'sd458715, 32'sd1683, 32'sd73465,
32'sd501347, 32'sd424870, 32'sd373017, 32'sd117086, 32'sd5651, 32'sd696479, 32'sd297176, 32'sd45610, 32'sd1236544, 32'sd905282,
32'sd750607, 32'sd205116, 32'sd109435, 32'sd412772, 32'sd318499, 32'sd147031, 32'sd568502, 32'sd25974, 32'sd23286, 32'sd897879,
32'sd118498, 32'sd103674, 32'sd725614, 32'sd372093, 32'sd324533, 32'sd315559, 32'sd162523, 32'sd191734, 32'sd51707, 32'sd593524,
32'sd52422, 32'sd665879, 32'sd49219, 32'sd39998, 32'sd144838, 32'sd572844, 32'sd336674, 32'sd236706, 32'sd190829, 32'sd362111,
32'sd7688, 32'sd124925, 32'sd855237, 32'sd69244, 32'sd191100, 32'sd292827, 32'sd168175, 32'sd55969, 32'sd199112, 32'sd200003,
32'sd3716, 32'sd333633, 32'sd366080, 32'sd45608, 32'sd254923, 32'sd162801, 32'sd4767, 32'sd38356, 32'sd249822, 32'sd102853,
32'sd15048, 32'sd451476, 32'sd81636, 32'sd1371218, 32'sd320676, 32'sd491883, 32'sd117951, 32'sd983307, 32'sd54138, 32'sd15733,
32'sd289062, 32'sd282044, 32'sd237750, 32'sd186740, 32'sd506836, 32'sd266470, 32'sd524105, 32'sd158713, 32'sd310581, 32'sd375956,
32'sd340962, 32'sd16964, 32'sd366188, 32'sd122247, 32'sd32392, 32'sd148660, 32'sd119272, 32'sd524415, 32'sd125085, 32'sd566453,
32'sd13875, 32'sd109644, 32'sd100614, 32'sd21761, 32'sd153114, 32'sd10906, 32'sd80547, 32'sd606181, 32'sd437738, 32'sd44781,
32'sd79902, 32'sd387229, 32'sd236527, 32'sd913252, 32'sd495765, 32'sd216386, 32'sd265420, 32'sd274516, 32'sd1012561, 32'sd48746,
32'sd346310, 32'sd317555, 32'sd300363, 32'sd563358, 32'sd258612, 32'sd277013, 32'sd536985, 32'sd85158, 32'sd207760, 32'sd18105,
32'sd288637, 32'sd730808, 32'sd56007, 32'sd2151, 32'sd269895, 32'sd69556, 32'sd10392, 32'sd43073, 32'sd73431, 32'sd52954,
32'sd6304, 32'sd300330, 32'sd340127, 32'sd476878, 32'sd247328, 32'sd358112, 32'sd17263, 32'sd353081, 32'sd1057471, 32'sd48168,
32'sd377607, 32'sd132859, 32'sd85236, 32'sd58194, 32'sd145805, 32'sd219224, 32'sd127120, 32'sd926271, 32'sd450354, 32'sd604195,
32'sd53256, 32'sd35276, 32'sd519770, 32'sd116254, 32'sd559287, 32'sd144659, 32'sd164444, 32'sd38908, 32'sd268417, 32'sd117652,
32'sd156848, 32'sd1909, 32'sd129378, 32'sd177638, 32'sd53967, 32'sd19121, 32'sd466199, 32'sd749885, 32'sd1093922, 32'sd38782,
32'sd54454, 32'sd75362, 32'sd33462, 32'sd201487, 32'sd20123, 32'sd203569, 32'sd212718, 32'sd168644, 32'sd409193, 32'sd851403,
32'sd158793, 32'sd713278, 32'sd368223, 32'sd108254, 32'sd196794, 32'sd793581, 32'sd380184, 32'sd884428, 32'sd677061, 32'sd219619,
32'sd136992, 32'sd31761, 32'sd353865, 32'sd40957, 32'sd16124, 32'sd231515, 32'sd22667, 32'sd263718, 32'sd333200, 32'sd236990,
32'sd135676, 32'sd380212, 32'sd17958, 32'sd672039, 32'sd192516, 32'sd12664, 32'sd42203, 32'sd324252, 32'sd280689, 32'sd49345,
32'sd859807, 32'sd35690, 32'sd139954, 32'sd855947, 32'sd502494, 32'sd337362, 32'sd283616, 32'sd292472, 32'sd44385, 32'sd574007,
32'sd257885, 32'sd190082, 32'sd158403, 32'sd336894, 32'sd137455, 32'sd336515, 32'sd991856, 32'sd55886, 32'sd338083, 32'sd206691,
32'sd318552, 32'sd194668, 32'sd240173, 32'sd129474, 32'sd422332, 32'sd6786, 32'sd175496, 32'sd16403, 32'sd151130, 32'sd936702,
32'sd510970, 32'sd265216, 32'sd89294, 32'sd568259, 32'sd22629, 32'sd122332, 32'sd52648, 32'sd42545, 32'sd5568, 32'sd336008,
32'sd705075, 32'sd174176, 32'sd134715, 32'sd41576, 32'sd48330, 32'sd583652, 32'sd150552, 32'sd414528, 32'sd131688, 32'sd683240,
32'sd260496, 32'sd2419, 32'sd36838, 32'sd74994, 32'sd219554, 32'sd195126, 32'sd36365, 32'sd404668, 32'sd65105, 32'sd98786,
32'sd301860, 32'sd351436, 32'sd142256, 32'sd560428, 32'sd422420, 32'sd961316, 32'sd154345, 32'sd165704, 32'sd243578, 32'sd151177,
32'sd113672, 32'sd440301, 32'sd108437, 32'sd144968, 32'sd415647, 32'sd304729, 32'sd117270, 32'sd269730, 32'sd15894, 32'sd63792,
32'sd245337, 32'sd172504, 32'sd71741, 32'sd141877, 32'sd367744, 32'sd139420, 32'sd620485, 32'sd345930, 32'sd41209, 32'sd394028,
32'sd444250, 32'sd196708, 32'sd299588, 32'sd90837, 32'sd372870, 32'sd181302, 32'sd77515, 32'sd125320, 32'sd186951, 32'sd144013,
32'sd141186, 32'sd96484, 32'sd132080, 32'sd8266, 32'sd260688, 32'sd182099, 32'sd238439, 32'sd506499, 32'sd289730, 32'sd166326,
32'sd121151, 32'sd164386, 32'sd146295, 32'sd388676, 32'sd566968, 32'sd102099, 32'sd233384, 32'sd363264, 32'sd341733, 32'sd12969,
32'sd244988, 32'sd389419, 32'sd160779, 32'sd478081, 32'sd376803, 32'sd154983, 32'sd123068, 32'sd894372, 32'sd1021315, 32'sd343607,
32'sd677019, 32'sd287930, 32'sd260022, 32'sd716328, 32'sd607454, 32'sd636437, 32'sd391014, 32'sd165165, 32'sd131820, 32'sd40153,
32'sd238603, 32'sd101348, 32'sd3387, 32'sd840933, 32'sd777911, 32'sd377181, 32'sd911521, 32'sd162015, 32'sd65048, 32'sd502834,
32'sd289002, 32'sd235458, 32'sd71756, 32'sd146344, 32'sd108779, 32'sd205603, 32'sd320079, 32'sd593697, 32'sd202971, 32'sd232575,
32'sd114464, 32'sd137715, 32'sd25925, 32'sd323034, 32'sd97944, 32'sd40055, 32'sd191418, 32'sd412449, 32'sd446719, 32'sd568813,
32'sd465628, 32'sd344814, 32'sd260938, 32'sd55481, 32'sd8415, 32'sd9250, 32'sd197932, 32'sd272299, 32'sd603018, 32'sd782297,
32'sd123549, 32'sd157371, 32'sd280937, 32'sd669733, 32'sd153219, 32'sd233607, 32'sd276837, 32'sd157052, 32'sd490842, 32'sd337175,
32'sd330644, 32'sd25428, 32'sd32153, 32'sd17524, 32'sd132513, 32'sd161903, 32'sd205680, 32'sd258475, 32'sd136872, 32'sd381612,
32'sd214128, 32'sd118411, 32'sd3722, 32'sd855142, 32'sd398031, 32'sd8742, 32'sd345120, 32'sd133625, 32'sd743166, 32'sd228842,
32'sd5224, 32'sd216654, 32'sd76654, 32'sd160709, 32'sd208138, 32'sd448708, 32'sd265451, 32'sd124680, 32'sd38608, 32'sd62133,
32'sd52946, 32'sd265930, 32'sd405128, 32'sd547202, 32'sd95109, 32'sd536727, 32'sd586628, 32'sd245652, 32'sd403120, 32'sd479307,
32'sd80816, 32'sd41532, 32'sd143706, 32'sd43121, 32'sd261390, 32'sd89141, 32'sd184393, 32'sd152192, 32'sd310417, 32'sd314611,
32'sd333011, 32'sd519339, 32'sd316410, 32'sd177805, 32'sd144657, 32'sd327138, 32'sd184631, 32'sd67295, 32'sd785584, 32'sd58580,
32'sd307560, 32'sd287562, 32'sd197370, 32'sd542238, 32'sd971944, 32'sd136102, 32'sd162186, 32'sd258388, 32'sd252227, 32'sd66382,
32'sd72259, 32'sd4335, 32'sd110935, 32'sd721687, 32'sd49332, 32'sd800850, 32'sd146987, 32'sd7888, 32'sd650016, 32'sd214536,
32'sd14844, 32'sd679007, 32'sd30009, 32'sd370072, 32'sd355499, 32'sd82687, 32'sd113013, 32'sd197697, 32'sd324594, 32'sd399900,
32'sd211550, 32'sd349726, 32'sd63633, 32'sd937574, 32'sd413700, 32'sd234391, 32'sd438554, 32'sd453564, 32'sd256727, 32'sd27758,
32'sd439282, 32'sd128993, 32'sd70486, 32'sd51298, 32'sd11702, 32'sd117823, 32'sd41287, 32'sd132591, 32'sd28079, 32'sd580318,
32'sd497760, 32'sd560497, 32'sd598474, 32'sd34852, 32'sd419257, 32'sd14423, 32'sd589029, 32'sd406243, 32'sd266749, 32'sd803303,
32'sd42601, 32'sd291232, 32'sd138696, 32'sd181074, 32'sd166164, 32'sd216613, 32'sd423514, 32'sd251291, 32'sd641470, 32'sd511465,
32'sd86783, 32'sd34099, 32'sd11922, 32'sd43126, 32'sd343679, 32'sd92567, 32'sd147684, 32'sd409217, 32'sd262594, 32'sd501064,
32'sd158859, 32'sd20894, 32'sd467960, 32'sd94252, 32'sd208342, 32'sd217403, 32'sd647802, 32'sd11682, 32'sd474295, 32'sd810931,
32'sd730117, 32'sd251836, 32'sd48292, 32'sd275237, 32'sd323409, 32'sd149593, 32'sd10501, 32'sd733497, 32'sd615956, 32'sd50730,
32'sd119625, 32'sd904722, 32'sd25580, 32'sd626849, 32'sd209799, 32'sd114928, 32'sd254715, 32'sd454433, 32'sd653075, 32'sd246493,
32'sd11213, 32'sd407833, 32'sd26343, 32'sd662328, 32'sd248248, 32'sd88220, 32'sd632727, 32'sd7492, 32'sd243348, 32'sd681,
32'sd19700, 32'sd916557, 32'sd248520, 32'sd281265, 32'sd319061, 32'sd131707, 32'sd17694, 32'sd126192, 32'sd561853, 32'sd53893,
32'sd968752, 32'sd1243252, 32'sd173655, 32'sd410800, 32'sd421676, 32'sd1053220, 32'sd237374, 32'sd279541, 32'sd290032, 32'sd10815,
32'sd1216518, 32'sd298158, 32'sd79596, 32'sd330074, 32'sd121849, 32'sd133354, 32'sd444202, 32'sd120223, 32'sd103418, 32'sd184858,
32'sd208077, 32'sd14564, 32'sd462057, 32'sd236590, 32'sd8804, 32'sd73277, 32'sd205196, 32'sd260882, 32'sd183014, 32'sd593114,
32'sd233749, 32'sd115747, 32'sd20156, 32'sd321010, 32'sd67424, 32'sd867304, 32'sd278593, 32'sd75963, 32'sd129198, 32'sd136543,
32'sd356096, 32'sd729848, 32'sd264134, 32'sd79688, 32'sd134534, 32'sd572633, 32'sd159876, 32'sd10335, 32'sd153709, 32'sd54112,
32'sd65356, 32'sd82744, 32'sd489332, 32'sd199494, 32'sd365130, 32'sd141642, 32'sd267549, 32'sd539221, 32'sd559237, 32'sd8842,
32'sd280438, 32'sd81342, 32'sd69280, 32'sd113511, 32'sd457321, 32'sd917309, 32'sd19334, 32'sd855771, 32'sd198405, 32'sd625789,
32'sd336261, 32'sd175641, 32'sd262426, 32'sd89040, 32'sd123727, 32'sd420460, 32'sd292468, 32'sd776690, 32'sd361962, 32'sd163373,
32'sd354833, 32'sd123045, 32'sd4776, 32'sd175780, 32'sd124008, 32'sd194661, 32'sd239243, 32'sd19669, 32'sd309258, 32'sd60346,
32'sd79031, 32'sd48488, 32'sd57050, 32'sd504347, 32'sd150481, 32'sd260923, 32'sd255646, 32'sd64966, 32'sd85608, 32'sd75788,
32'sd36830, 32'sd603032, 32'sd5980, 32'sd102207, 32'sd82096, 32'sd119741, 32'sd52705, 32'sd84303, 32'sd169320, 32'sd73297,
32'sd119678, 32'sd313905, 32'sd268853, 32'sd89382, 32'sd150011, 32'sd362285, 32'sd133708, 32'sd381836, 32'sd41868, 32'sd77100,
32'sd231454, 32'sd6182, 32'sd345303, 32'sd468286, 32'sd706841, 32'sd817, 32'sd22560, 32'sd44724, 32'sd166572, 32'sd85642,
32'sd5496, 32'sd174737, 32'sd276354, 32'sd198648, 32'sd373823, 32'sd440378, 32'sd317430, 32'sd405449, 32'sd239904, 32'sd227563,
32'sd155626, 32'sd142215, 32'sd101472, 32'sd119820, 32'sd29587, 32'sd179109, 32'sd450750, 32'sd66529, 32'sd68943, 32'sd191623,
32'sd26453, 32'sd204114, 32'sd76077, 32'sd66131, 32'sd110232, 32'sd360412, 32'sd225434, 32'sd644446, 32'sd150224, 32'sd712898,
32'sd43823, 32'sd175510, 32'sd44706, 32'sd746757, 32'sd156176, 32'sd121107, 32'sd1357, 32'sd309333, 32'sd43937, 32'sd138335,
32'sd300539, 32'sd40063, 32'sd250074, 32'sd739253, 32'sd105448, 32'sd539400, 32'sd205757, 32'sd844899, 32'sd19945, 32'sd999514,
32'sd80936, 32'sd17707, 32'sd47441, 32'sd21264, 32'sd124184, 32'sd133877, 32'sd317620, 32'sd33711, 32'sd236973, 32'sd18235,
32'sd108610, 32'sd66482, 32'sd96828, 32'sd45085, 32'sd501149, 32'sd467078, 32'sd10413, 32'sd317764, 32'sd68818, 32'sd594402,
32'sd440832, 32'sd139499, 32'sd50214, 32'sd264247, 32'sd57360, 32'sd453685, 32'sd235880, 32'sd153750, 32'sd39320, 32'sd187746,
32'sd10548, 32'sd536322, 32'sd177582, 32'sd361664, 32'sd337094, 32'sd191780, 32'sd610635, 32'sd306863, 32'sd377013, 32'sd92148,
32'sd104373, 32'sd113117, 32'sd260773, 32'sd546445, 32'sd597801, 32'sd50713, 32'sd48601, 32'sd376546, 32'sd561274, 32'sd1869,
32'sd48315, 32'sd98829, 32'sd434747, 32'sd176082, 32'sd182293, 32'sd31257, 32'sd373488, 32'sd386436, 32'sd139885, 32'sd152104,
32'sd358198, 32'sd371376, 32'sd170255, 32'sd17430, 32'sd238990, 32'sd473395, 32'sd232770, 32'sd499005, 32'sd1211076, 32'sd246892,
32'sd812018, 32'sd859311, 32'sd64951, 32'sd259440, 32'sd76832, 32'sd10203, 32'sd705765, 32'sd414088, 32'sd271523, 32'sd235144,
32'sd409921, 32'sd101785, 32'sd87325, 32'sd392752, 32'sd28821, 32'sd141877, 32'sd668374, 32'sd75412, 32'sd349222, 32'sd132854,
32'sd286533, 32'sd339155, 32'sd356698, 32'sd55611, 32'sd21791, 32'sd1019961, 32'sd83394, 32'sd78338, 32'sd277918, 32'sd102083,
32'sd600113, 32'sd105073, 32'sd609915, 32'sd109745, 32'sd64836, 32'sd193972, 32'sd377055, 32'sd386910, 32'sd73834, 32'sd71717,
32'sd288410, 32'sd71762, 32'sd119066, 32'sd26953, 32'sd4250, 32'sd106368, 32'sd135741, 32'sd60171, 32'sd134417, 32'sd52693,
32'sd196335, 32'sd135516, 32'sd165488, 32'sd874624, 32'sd52992, 32'sd8928, 32'sd238160, 32'sd183767, 32'sd85959, 32'sd208702,
32'sd47283, 32'sd271604, 32'sd29231, 32'sd30171, 32'sd280527, 32'sd773620, 32'sd126735, 32'sd21829, 32'sd110764, 32'sd305926,
32'sd86391, 32'sd35001, 32'sd629709, 32'sd321762, 32'sd81417, 32'sd288472, 32'sd157381, 32'sd129627, 32'sd127018, 32'sd621457,
32'sd57920, 32'sd164694, 32'sd174336, 32'sd137474, 32'sd140814, 32'sd556237, 32'sd439, 32'sd205427, 32'sd340488, 32'sd240444,
32'sd183279, 32'sd108620, 32'sd76952, 32'sd690169, 32'sd103157, 32'sd130862, 32'sd54839, 32'sd14963, 32'sd562258, 32'sd156935,
32'sd717217, 32'sd879586, 32'sd410408, 32'sd8221, 32'sd413101, 32'sd1057193, 32'sd564462, 32'sd336348, 32'sd160795, 32'sd228359,
32'sd686985, 32'sd4758, 32'sd261070, 32'sd495711, 32'sd432887, 32'sd112673, 32'sd156800, 32'sd142792, 32'sd159240, 32'sd18811,
32'sd87666, 32'sd227238, 32'sd160114, 32'sd195495, 32'sd198415, 32'sd106516, 32'sd550569, 32'sd250232, 32'sd730772, 32'sd359017,
32'sd130702, 32'sd13575, 32'sd146236, 32'sd499753, 32'sd371424, 32'sd889709, 32'sd120695, 32'sd71036, 32'sd216008, 32'sd814276,
32'sd178094, 32'sd159097, 32'sd308139, 32'sd221246, 32'sd369679, 32'sd1176, 32'sd45163, 32'sd639377, 32'sd218133, 32'sd82694,
32'sd394473, 32'sd260888, 32'sd69866, 32'sd331719, 32'sd48992, 32'sd417961, 32'sd189720, 32'sd197676, 32'sd63142, 32'sd443441,
32'sd218996, 32'sd478552, 32'sd449412, 32'sd593002, 32'sd749306, 32'sd612446, 32'sd188877, 32'sd745057, 32'sd82937, 32'sd549680,
32'sd89577, 32'sd89051, 32'sd249882, 32'sd19637, 32'sd381820, 32'sd286360, 32'sd36876, 32'sd116794, 32'sd48755, 32'sd175630,
32'sd251486, 32'sd88960, 32'sd247823, 32'sd206730, 32'sd490494, 32'sd140634, 32'sd480118, 32'sd225059, 32'sd291484, 32'sd204860,
32'sd546879, 32'sd168528, 32'sd423760, 32'sd69434, 32'sd152866, 32'sd336969, 32'sd70268, 32'sd47988, 32'sd40987, 32'sd84875,
32'sd303160, 32'sd814656, 32'sd276988, 32'sd55195, 32'sd848812, 32'sd144960, 32'sd126547, 32'sd98047, 32'sd233636, 32'sd484854,
32'sd115720, 32'sd528369, 32'sd409780, 32'sd123420, 32'sd51128, 32'sd194876, 32'sd190285, 32'sd225579, 32'sd121238, 32'sd218160,
32'sd585632, 32'sd2475, 32'sd68478, 32'sd165104, 32'sd522290, 32'sd120417, 32'sd308443, 32'sd90008, 32'sd241605, 32'sd255619,
32'sd980891, 32'sd328199, 32'sd100352, 32'sd89292, 32'sd3486, 32'sd172938, 32'sd7649, 32'sd751, 32'sd199436, 32'sd338098,
32'sd4255, 32'sd162016, 32'sd403070, 32'sd503649, 32'sd120305, 32'sd173625, 32'sd30540, 32'sd784775, 32'sd411247, 32'sd213991,
32'sd259272, 32'sd363454, 32'sd123237, 32'sd166898, 32'sd780672, 32'sd45521, 32'sd361368, 32'sd694747, 32'sd139542, 32'sd1800,
32'sd15404, 32'sd34889, 32'sd146331, 32'sd44640, 32'sd85841, 32'sd1086352, 32'sd289757, 32'sd29622, 32'sd143948, 32'sd1613389,
32'sd292927, 32'sd344124, 32'sd286538, 32'sd454947, 32'sd678848, 32'sd345379, 32'sd34139, 32'sd1113430, 32'sd303353, 32'sd114163,
32'sd321466, 32'sd367667, 32'sd117150, 32'sd28899, 32'sd673598, 32'sd155239, 32'sd665836, 32'sd201512, 32'sd255481, 32'sd82181,
32'sd466431, 32'sd177756, 32'sd370896, 32'sd157793, 32'sd512977, 32'sd50948, 32'sd431690, 32'sd31297, 32'sd793129, 32'sd31754,
32'sd286035, 32'sd149731, 32'sd580017, 32'sd254955, 32'sd487892, 32'sd591684, 32'sd1381999, 32'sd210494, 32'sd5841, 32'sd665355,
32'sd296822, 32'sd428370, 32'sd93823, 32'sd445648, 32'sd338626, 32'sd238455, 32'sd400557, 32'sd87328, 32'sd310808, 32'sd982611,
32'sd171753, 32'sd477029, 32'sd473753, 32'sd332898, 32'sd62687, 32'sd453861, 32'sd54756, 32'sd91885, 32'sd665957, 32'sd125652,
32'sd39245, 32'sd23790, 32'sd232682, 32'sd80115, 32'sd220540, 32'sd113669, 32'sd432489, 32'sd81150, 32'sd304812, 32'sd92168,
32'sd235406, 32'sd315050, 32'sd44099, 32'sd676279, 32'sd94390, 32'sd670747, 32'sd204314, 32'sd459418, 32'sd6300, 32'sd297542,
32'sd168224, 32'sd911665, 32'sd1065790, 32'sd220165, 32'sd472014, 32'sd134792, 32'sd15099, 32'sd87536, 32'sd804394, 32'sd306535,
32'sd484148, 32'sd52901, 32'sd90376, 32'sd19116, 32'sd309597, 32'sd170818, 32'sd13170, 32'sd150358, 32'sd178671, 32'sd128296,
32'sd152544, 32'sd135454, 32'sd476203, 32'sd34423, 32'sd75148, 32'sd513960, 32'sd87239, 32'sd29448, 32'sd183545, 32'sd82631,
32'sd428208, 32'sd109250, 32'sd222229, 32'sd76103, 32'sd643753, 32'sd193653, 32'sd354774, 32'sd696352, 32'sd62373, 32'sd18889,
32'sd297344, 32'sd270326, 32'sd168091, 32'sd154167, 32'sd51052, 32'sd231785, 32'sd295704, 32'sd255902, 32'sd290915, 32'sd382195,
32'sd87035, 32'sd58233, 32'sd449920, 32'sd203705, 32'sd80706, 32'sd742086, 32'sd630195, 32'sd166970, 32'sd71649, 32'sd218002,
32'sd107638, 32'sd34213, 32'sd291343, 32'sd263085, 32'sd6901, 32'sd47839, 32'sd302463, 32'sd213154, 32'sd94459, 32'sd172221,
32'sd47791, 32'sd116240, 32'sd177955, 32'sd898936, 32'sd423603, 32'sd197504, 32'sd204491, 32'sd157289, 32'sd701575, 32'sd146123,
32'sd439285, 32'sd489784, 32'sd21910, 32'sd57303, 32'sd94884, 32'sd187184, 32'sd50422, 32'sd105690, 32'sd110752, 32'sd162035,
32'sd830280, 32'sd400561, 32'sd365357, 32'sd403531, 32'sd695564, 32'sd138572, 32'sd150343, 32'sd358207, 32'sd975569, 32'sd715776,
32'sd277008, 32'sd626489, 32'sd118733, 32'sd466566, 32'sd26009, 32'sd225980, 32'sd57808, 32'sd242525, 32'sd477001, 32'sd113756,
32'sd227702, 32'sd286472, 32'sd955700, 32'sd122721, 32'sd534424, 32'sd817369, 32'sd18522, 32'sd32038, 32'sd107546, 32'sd363468,
32'sd222434, 32'sd292236, 32'sd459434, 32'sd242347, 32'sd243460, 32'sd257979, 32'sd231402, 32'sd485717, 32'sd262803, 32'sd645701,
32'sd169293, 32'sd832635, 32'sd266710, 32'sd244604, 32'sd3552, 32'sd39977, 32'sd226596, 32'sd252048, 32'sd4544, 32'sd77071,
32'sd319203, 32'sd90045, 32'sd1028157, 32'sd426835, 32'sd141337, 32'sd377620, 32'sd25977, 32'sd99365, 32'sd36403, 32'sd156667,
32'sd24428, 32'sd143141, 32'sd768785, 32'sd297280, 32'sd381040, 32'sd241851, 32'sd274111, 32'sd411625, 32'sd486454, 32'sd13254,
32'sd96790, 32'sd171768, 32'sd61950, 32'sd321984, 32'sd321007, 32'sd170329, 32'sd191730, 32'sd182907, 32'sd866264, 32'sd383854,
32'sd213281, 32'sd57782, 32'sd384828, 32'sd78398, 32'sd643198, 32'sd12157, 32'sd1220751, 32'sd180864, 32'sd6639, 32'sd129358,
32'sd63598, 32'sd93979, 32'sd56626, 32'sd271013, 32'sd19004, 32'sd141302, 32'sd371869, 32'sd49423, 32'sd462919, 32'sd164813,
32'sd112152, 32'sd388470, 32'sd254981, 32'sd42010, 32'sd66416, 32'sd142071, 32'sd15022, 32'sd383764, 32'sd109325, 32'sd199998,
32'sd331393, 32'sd353245, 32'sd312534, 32'sd179057, 32'sd282338, 32'sd283555, 32'sd745647, 32'sd328828, 32'sd257450, 32'sd19705,
32'sd430312, 32'sd18779, 32'sd30188, 32'sd498582, 32'sd214029, 32'sd15381, 32'sd86273, 32'sd101736, 32'sd274645, 32'sd77952,
32'sd454748, 32'sd361568, 32'sd363654, 32'sd85193, 32'sd30112, 32'sd183890, 32'sd8349, 32'sd63175, 32'sd793507, 32'sd112405,
32'sd107697, 32'sd98578, 32'sd153185, 32'sd512122, 32'sd154156, 32'sd146880, 32'sd66435, 32'sd423489, 32'sd80022, 32'sd68408,
32'sd336324, 32'sd6152, 32'sd1739, 32'sd543013, 32'sd857458, 32'sd45143, 32'sd472382, 32'sd130839, 32'sd273856, 32'sd820682,
32'sd7642, 32'sd151015, 32'sd812018, 32'sd93419, 32'sd75968, 32'sd42680, 32'sd41382, 32'sd146264, 32'sd155645, 32'sd542331,
32'sd126509, 32'sd231222, 32'sd854703, 32'sd12852, 32'sd239883, 32'sd314163, 32'sd33597, 32'sd178493, 32'sd34217, 32'sd515415,
32'sd69505, 32'sd529440, 32'sd71764, 32'sd156261, 32'sd134750, 32'sd622167, 32'sd374965, 32'sd470147, 32'sd3394, 32'sd36580,
32'sd280621, 32'sd67858, 32'sd19226, 32'sd139484, 32'sd977184, 32'sd251762, 32'sd590230, 32'sd391236, 32'sd207348, 32'sd857376,
32'sd14575, 32'sd150273, 32'sd470, 32'sd150016, 32'sd49179, 32'sd78388, 32'sd306346, 32'sd8226, 32'sd409394, 32'sd204893,
32'sd592091, 32'sd241125, 32'sd94076, 32'sd112052, 32'sd100102, 32'sd531049, 32'sd632753, 32'sd431622, 32'sd603356, 32'sd523129,
32'sd557181, 32'sd840287, 32'sd12592, 32'sd302246, 32'sd107024, 32'sd508196, 32'sd18694, 32'sd51957, 32'sd465764, 32'sd493599,
32'sd351958, 32'sd187134, 32'sd377184, 32'sd652462, 32'sd86232, 32'sd329548, 32'sd374718, 32'sd314738, 32'sd170472, 32'sd695026,
32'sd165290, 32'sd14617, 32'sd335677, 32'sd14956, 32'sd170011, 32'sd72042, 32'sd4598, 32'sd107496, 32'sd153907, 32'sd935307,
32'sd56253, 32'sd162818, 32'sd441269, 32'sd659206, 32'sd59942, 32'sd120003, 32'sd105930, 32'sd720003, 32'sd241749, 32'sd266244,
32'sd178900, 32'sd298318, 32'sd229430, 32'sd145210, 32'sd109692, 32'sd42521, 32'sd94579, 32'sd254591, 32'sd281588, 32'sd240483,
32'sd220061, 32'sd114750, 32'sd6526, 32'sd20357, 32'sd243156, 32'sd488865, 32'sd104752, 32'sd242235, 32'sd478632, 32'sd163942,
32'sd967865, 32'sd134880, 32'sd121227, 32'sd190951, 32'sd370005, 32'sd165606, 32'sd992, 32'sd66525, 32'sd669659, 32'sd16692,
32'sd15517, 32'sd157176, 32'sd122788, 32'sd55820, 32'sd146965, 32'sd276604, 32'sd39411, 32'sd341729, 32'sd62382, 32'sd14043,
32'sd688678, 32'sd603255, 32'sd385978, 32'sd212533, 32'sd771804, 32'sd279675, 32'sd514663, 32'sd302685, 32'sd473722, 32'sd96866,
32'sd32380, 32'sd416492, 32'sd652216, 32'sd150989, 32'sd127653, 32'sd1836, 32'sd24601, 32'sd283999, 32'sd30658, 32'sd416862,
32'sd208602, 32'sd92065, 32'sd293166, 32'sd203673, 32'sd276414, 32'sd136909, 32'sd251678, 32'sd32415, 32'sd73779, 32'sd20471,
32'sd6912, 32'sd112756, 32'sd97772, 32'sd351536, 32'sd25662, 32'sd177150, 32'sd144537, 32'sd461691, 32'sd95421, 32'sd359039,
32'sd7798, 32'sd3290, 32'sd46475, 32'sd273677, 32'sd72010, 32'sd159897, 32'sd7296, 32'sd70149, 32'sd310348, 32'sd114140,
32'sd504644, 32'sd427373, 32'sd729919, 32'sd454058, 32'sd275807, 32'sd181111, 32'sd764620, 32'sd192160, 32'sd76846, 32'sd220900,
32'sd345004, 32'sd218523, 32'sd542428, 32'sd64897, 32'sd234380, 32'sd457626, 32'sd141098, 32'sd69218, 32'sd36616, 32'sd28929,
32'sd287264, 32'sd506789, 32'sd887080, 32'sd277194, 32'sd218883, 32'sd93039, 32'sd101934, 32'sd301258, 32'sd288892, 32'sd523652,
32'sd575164, 32'sd803809, 32'sd129629, 32'sd236160, 32'sd183382, 32'sd7830, 32'sd93265, 32'sd250734, 32'sd46546, 32'sd600210,
32'sd501313, 32'sd109884, 32'sd425610, 32'sd317501, 32'sd268197, 32'sd241732, 32'sd607987, 32'sd205896, 32'sd6815, 32'sd10895,
32'sd64541, 32'sd158582, 32'sd332199, 32'sd551370, 32'sd719358, 32'sd656971, 32'sd118050, 32'sd55829, 32'sd111440, 32'sd22860,
32'sd68519, 32'sd445514, 32'sd330441, 32'sd52469, 32'sd233416, 32'sd188865, 32'sd461509, 32'sd645195, 32'sd193479, 32'sd203165,
32'sd209910, 32'sd202823, 32'sd496515, 32'sd618065, 32'sd479750, 32'sd289452, 32'sd301794, 32'sd83110, 32'sd10436, 32'sd36839,
32'sd23865, 32'sd196215, 32'sd292338, 32'sd40080, 32'sd2384, 32'sd109240, 32'sd1901, 32'sd632161, 32'sd654100, 32'sd11771,
32'sd142107, 32'sd12289, 32'sd540193, 32'sd98551, 32'sd379148, 32'sd304462, 32'sd433922, 32'sd405842, 32'sd333292, 32'sd35838,
32'sd148359, 32'sd32166, 32'sd381923, 32'sd106240, 32'sd30367, 32'sd114578, 32'sd878696, 32'sd340233, 32'sd130869, 32'sd206124,
32'sd341537, 32'sd82772, 32'sd54327, 32'sd516698, 32'sd592643, 32'sd405307, 32'sd99250, 32'sd326150, 32'sd17746, 32'sd6867,
32'sd81985, 32'sd558374, 32'sd370803, 32'sd403149, 32'sd183924, 32'sd353481, 32'sd767912, 32'sd294429, 32'sd370719, 32'sd342783,
32'sd363803, 32'sd658724, 32'sd629058, 32'sd119818, 32'sd210321, 32'sd242710, 32'sd250827, 32'sd370650, 32'sd108512, 32'sd70340,
32'sd136522, 32'sd184463, 32'sd34132, 32'sd395465, 32'sd173209, 32'sd416579, 32'sd114926, 32'sd454905, 32'sd77745, 32'sd423448,
32'sd119638, 32'sd305092, 32'sd62886, 32'sd290608, 32'sd101368, 32'sd514038, 32'sd372124, 32'sd368316, 32'sd117743, 32'sd322121,
32'sd101451, 32'sd20751, 32'sd238641, 32'sd498782, 32'sd110529, 32'sd123221, 32'sd643215, 32'sd35052, 32'sd27788, 32'sd321770,
32'sd620173, 32'sd206130, 32'sd155552, 32'sd30171, 32'sd254406, 32'sd671447, 32'sd408378, 32'sd21874, 32'sd33374, 32'sd203881,
32'sd149146, 32'sd702515, 32'sd203763, 32'sd297921, 32'sd130371, 32'sd22346, 32'sd329059, 32'sd309302, 32'sd74763, 32'sd302662,
32'sd393688, 32'sd93438, 32'sd384998, 32'sd131248, 32'sd57116, 32'sd309442, 32'sd69463, 32'sd7723, 32'sd468620, 32'sd90500,
32'sd190268, 32'sd79080, 32'sd82612, 32'sd796929, 32'sd161861, 32'sd707115, 32'sd201004, 32'sd102951, 32'sd250931, 32'sd24498,
32'sd243571, 32'sd52199, 32'sd42664, 32'sd397071, 32'sd681534, 32'sd395846, 32'sd373158, 32'sd7238, 32'sd111904, 32'sd297996,
32'sd181142, 32'sd364126, 32'sd493364, 32'sd633034, 32'sd188071, 32'sd175129, 32'sd90455, 32'sd106612, 32'sd116023, 32'sd106039,
32'sd119546, 32'sd166482, 32'sd148669, 32'sd173662, 32'sd189974, 32'sd78909, 32'sd588772, 32'sd159183, 32'sd808878, 32'sd146979,
32'sd86155, 32'sd284628, 32'sd146947, 32'sd105689, 32'sd734710, 32'sd394192, 32'sd59711, 32'sd64169, 32'sd911493, 32'sd712454,
32'sd381161, 32'sd689909, 32'sd18289, 32'sd107740, 32'sd92901, 32'sd176224, 32'sd78041, 32'sd133, 32'sd66394, 32'sd225219,
32'sd88139, 32'sd502972, 32'sd7354, 32'sd29419, 32'sd26732, 32'sd291447, 32'sd99069, 32'sd121815, 32'sd100458, 32'sd375164,
32'sd37361, 32'sd178160, 32'sd89309, 32'sd345019, 32'sd202812, 32'sd301023, 32'sd426360, 32'sd24330, 32'sd604662, 32'sd245395,
32'sd262900, 32'sd184993, 32'sd1087265, 32'sd779270, 32'sd525807, 32'sd558541, 32'sd40, 32'sd346293, 32'sd36750, 32'sd262050,
32'sd322392, 32'sd25922, 32'sd406395, 32'sd508896, 32'sd413116, 32'sd119837, 32'sd3659, 32'sd583430, 32'sd125586, 32'sd275825,
32'sd174397, 32'sd252998, 32'sd566660, 32'sd766722, 32'sd350984, 32'sd290070, 32'sd62918, 32'sd148680, 32'sd248044, 32'sd50597,
32'sd163898, 32'sd283579, 32'sd9165, 32'sd14479, 32'sd134816, 32'sd109760, 32'sd620480, 32'sd488634, 32'sd1030577, 32'sd115766,
32'sd209355, 32'sd99237, 32'sd48297, 32'sd40678, 32'sd96151, 32'sd339269, 32'sd869448, 32'sd696202, 32'sd458770, 32'sd632681,
32'sd848286, 32'sd69217, 32'sd249109, 32'sd437027, 32'sd122165, 32'sd229052, 32'sd480858, 32'sd72284, 32'sd172099, 32'sd25129,
32'sd761192, 32'sd57867, 32'sd177251, 32'sd565869, 32'sd300340, 32'sd341726, 32'sd64698, 32'sd139629, 32'sd96559, 32'sd130846,
32'sd309810, 32'sd229921, 32'sd381880, 32'sd211722, 32'sd102459, 32'sd400565, 32'sd15598, 32'sd24642, 32'sd157405, 32'sd191685,
32'sd16268, 32'sd495736, 32'sd32525, 32'sd58605, 32'sd308863, 32'sd414578, 32'sd208402, 32'sd116512, 32'sd147383, 32'sd43438,
32'sd455586, 32'sd244773, 32'sd174748, 32'sd461436, 32'sd276357, 32'sd153879, 32'sd578934, 32'sd511640, 32'sd408591, 32'sd185192,
32'sd146752, 32'sd194700, 32'sd35988, 32'sd395160, 32'sd36168, 32'sd747990, 32'sd407073, 32'sd99602, 32'sd62176, 32'sd589186,
32'sd228101, 32'sd132581, 32'sd259761, 32'sd42878, 32'sd354705, 32'sd121092, 32'sd596441, 32'sd355706, 32'sd293640, 32'sd501253,
32'sd335427, 32'sd174234, 32'sd189749, 32'sd8096, 32'sd441576, 32'sd740005, 32'sd24242, 32'sd718648, 32'sd117486, 32'sd11225,
32'sd485232, 32'sd867146, 32'sd527286, 32'sd23988, 32'sd64002, 32'sd129893, 32'sd940752, 32'sd172355, 32'sd84724, 32'sd626837,
32'sd428917, 32'sd578809, 32'sd372763, 32'sd126084, 32'sd214214, 32'sd66272, 32'sd37739, 32'sd303004, 32'sd26842, 32'sd110370,
32'sd409988, 32'sd13452, 32'sd34242, 32'sd855895, 32'sd219902, 32'sd8204, 32'sd16289, 32'sd438493, 32'sd61985, 32'sd497093,
32'sd297269, 32'sd77222, 32'sd337652, 32'sd12453, 32'sd311602, 32'sd512771, 32'sd421647, 32'sd77272, 32'sd279762, 32'sd5652,
32'sd78409, 32'sd79261, 32'sd159504, 32'sd1118984, 32'sd368280, 32'sd157738, 32'sd72879, 32'sd196073, 32'sd352830, 32'sd391563,
32'sd48206, 32'sd312655, 32'sd72344, 32'sd181590, 32'sd800812, 32'sd39076, 32'sd99132, 32'sd399313, 32'sd61296, 32'sd294897,
32'sd23374, 32'sd15142, 32'sd828284, 32'sd120901, 32'sd764475, 32'sd287775, 32'sd788592, 32'sd266331, 32'sd563874, 32'sd97501,
32'sd98690, 32'sd533250, 32'sd363686, 32'sd36027, 32'sd830466, 32'sd557863, 32'sd371948, 32'sd68373, 32'sd56552, 32'sd253125,
32'sd15278, 32'sd55648, 32'sd188178, 32'sd20672, 32'sd23868, 32'sd199636, 32'sd154846, 32'sd182955, 32'sd553305, 32'sd388797,
32'sd577786, 32'sd552835, 32'sd337087, 32'sd15193, 32'sd199729, 32'sd127310, 32'sd394122, 32'sd475320, 32'sd684012, 32'sd36347,
32'sd159458, 32'sd37224, 32'sd221955, 32'sd144031, 32'sd65698, 32'sd326869, 32'sd150295, 32'sd45492, 32'sd70105, 32'sd173968,
32'sd171235, 32'sd88309, 32'sd89999, 32'sd370477, 32'sd120106, 32'sd964427, 32'sd297461, 32'sd238200, 32'sd889470, 32'sd916174,
32'sd98930, 32'sd13882, 32'sd143418, 32'sd314348, 32'sd33203, 32'sd229427, 32'sd273900, 32'sd515889, 32'sd455260, 32'sd213537,
32'sd121894, 32'sd175830, 32'sd691100, 32'sd660422, 32'sd433068, 32'sd155459, 32'sd299346, 32'sd35864, 32'sd68706, 32'sd213369,
32'sd158659, 32'sd260240, 32'sd489785, 32'sd33630, 32'sd58612, 32'sd67630, 32'sd84655, 32'sd371685, 32'sd350872, 32'sd271034,
32'sd222704, 32'sd142892, 32'sd111823, 32'sd196368, 32'sd2269, 32'sd16713, 32'sd71010, 32'sd435934, 32'sd843128, 32'sd5934,
32'sd316457, 32'sd245654, 32'sd801752, 32'sd15309, 32'sd426846, 32'sd98200, 32'sd12866, 32'sd550258, 32'sd82120, 32'sd86828,
32'sd42486, 32'sd16580, 32'sd735224, 32'sd331043, 32'sd325501, 32'sd228244, 32'sd5589, 32'sd943683, 32'sd48706, 32'sd49496,
32'sd299363, 32'sd133400, 32'sd276537, 32'sd56104, 32'sd370167, 32'sd136741, 32'sd187974, 32'sd271288, 32'sd184172, 32'sd85662,
32'sd510655, 32'sd66839, 32'sd35305, 32'sd583222, 32'sd143690, 32'sd602863, 32'sd399730, 32'sd129706, 32'sd161415, 32'sd79705,
32'sd141864, 32'sd89162, 32'sd185551, 32'sd253239, 32'sd200212, 32'sd100667, 32'sd55205, 32'sd316999, 32'sd52747, 32'sd164298,
32'sd251221, 32'sd529539, 32'sd499385, 32'sd421870, 32'sd398402, 32'sd107566, 32'sd142521, 32'sd586044, 32'sd987966, 32'sd63124,
32'sd826429, 32'sd607440, 32'sd508393, 32'sd919630, 32'sd192996, 32'sd741864, 32'sd738183, 32'sd372878, 32'sd296964, 32'sd222884,
32'sd1153553, 32'sd106580, 32'sd21762, 32'sd396549, 32'sd163116, 32'sd63406, 32'sd180651, 32'sd52227, 32'sd296655, 32'sd243197,
32'sd628914, 32'sd107155, 32'sd86546, 32'sd263880, 32'sd761451, 32'sd894028, 32'sd58794, 32'sd206981, 32'sd94804, 32'sd331067,
32'sd259306, 32'sd144614, 32'sd4656, 32'sd210036, 32'sd196219, 32'sd190981, 32'sd329184, 32'sd18897, 32'sd802632, 32'sd268636,
32'sd155597, 32'sd106717, 32'sd123502, 32'sd47353, 32'sd93081, 32'sd163278, 32'sd218668, 32'sd674368, 32'sd224611, 32'sd345410,
32'sd306028, 32'sd174146, 32'sd718980, 32'sd215965, 32'sd235589, 32'sd109566, 32'sd636617, 32'sd741936, 32'sd54071, 32'sd168294,
32'sd539464, 32'sd16288, 32'sd135005, 32'sd426122, 32'sd185492, 32'sd143839, 32'sd285274, 32'sd540989, 32'sd344806, 32'sd359392,
32'sd136956, 32'sd555626, 32'sd84042, 32'sd100003, 32'sd157800, 32'sd308362, 32'sd160645, 32'sd562770, 32'sd155105, 32'sd191532,
32'sd340670, 32'sd79443, 32'sd495782, 32'sd878182, 32'sd10533, 32'sd1056949, 32'sd323967, 32'sd151190, 32'sd407938, 32'sd173953,
32'sd450604, 32'sd6469, 32'sd53679, 32'sd167920, 32'sd184823, 32'sd100837, 32'sd100784, 32'sd236804, 32'sd541384, 32'sd671268,
32'sd206476, 32'sd244488, 32'sd68344, 32'sd31986, 32'sd53511, 32'sd489164, 32'sd90106, 32'sd10612, 32'sd414087, 32'sd25370,
32'sd90256, 32'sd42945, 32'sd210572, 32'sd275064, 32'sd10434, 32'sd86696, 32'sd12956, 32'sd320051, 32'sd182702, 32'sd48373,
32'sd661001, 32'sd333254, 32'sd310646, 32'sd85450, 32'sd1095, 32'sd118232, 32'sd71966, 32'sd352077, 32'sd484768, 32'sd723168,
32'sd399366, 32'sd321286, 32'sd676678, 32'sd1274675, 32'sd12010, 32'sd181, 32'sd378647, 32'sd1175926, 32'sd202957, 32'sd183092,
32'sd330042, 32'sd449511, 32'sd281669, 32'sd61165, 32'sd14347, 32'sd177725, 32'sd128292, 32'sd541290, 32'sd110568, 32'sd1109039,
32'sd302760, 32'sd133593, 32'sd146564, 32'sd134045, 32'sd53068, 32'sd76832, 32'sd325178, 32'sd70571, 32'sd6792, 32'sd126463,
32'sd647146, 32'sd601789, 32'sd221814, 32'sd85290, 32'sd45838, 32'sd125622, 32'sd141040, 32'sd16252, 32'sd186299, 32'sd231863,
32'sd337962, 32'sd141909, 32'sd924574, 32'sd153405, 32'sd164072, 32'sd89940, 32'sd100118, 32'sd614414, 32'sd83828, 32'sd289216,
32'sd304462, 32'sd282428, 32'sd352565, 32'sd81654, 32'sd233409, 32'sd254660, 32'sd228919, 32'sd184660, 32'sd101011, 32'sd294193,
32'sd379472, 32'sd35730, 32'sd23353, 32'sd397119, 32'sd208454, 32'sd122497, 32'sd156173, 32'sd282068, 32'sd434671, 32'sd143548,
32'sd77238, 32'sd322823, 32'sd102039, 32'sd408996, 32'sd149810, 32'sd179166, 32'sd265399, 32'sd190450, 32'sd395597, 32'sd752839,
32'sd406759, 32'sd14952, 32'sd405138, 32'sd2794, 32'sd281634, 32'sd119958, 32'sd153611, 32'sd618646, 32'sd312861, 32'sd296656,
32'sd127922, 32'sd52188, 32'sd290606, 32'sd42208, 32'sd339216, 32'sd36951, 32'sd159811, 32'sd507948, 32'sd50829, 32'sd196115,
32'sd150859, 32'sd104470, 32'sd76318, 32'sd139982, 32'sd471853, 32'sd26518, 32'sd171522, 32'sd25357, 32'sd137334, 32'sd6408,
32'sd2541, 32'sd461415, 32'sd2837, 32'sd929235, 32'sd669303, 32'sd75705, 32'sd628805, 32'sd287622, 32'sd114967, 32'sd53802,
32'sd150215, 32'sd557457, 32'sd273416, 32'sd95666, 32'sd151397, 32'sd222740, 32'sd64041, 32'sd541891, 32'sd592516, 32'sd39487,
32'sd4747, 32'sd572552, 32'sd286310, 32'sd153000, 32'sd118671, 32'sd87707, 32'sd21654, 32'sd58971, 32'sd137861, 32'sd296824,
32'sd93182, 32'sd308157, 32'sd72103, 32'sd404618, 32'sd728066, 32'sd158207, 32'sd18143, 32'sd365649, 32'sd618023, 32'sd116589,
32'sd682032, 32'sd289298, 32'sd59271, 32'sd898119, 32'sd41986, 32'sd234507, 32'sd115528, 32'sd414001, 32'sd518276, 32'sd324472,
32'sd244264, 32'sd1032346, 32'sd635057, 32'sd18021, 32'sd170379, 32'sd135132, 32'sd116275, 32'sd322717, 32'sd11217, 32'sd511010,
32'sd370442, 32'sd408621, 32'sd31730, 32'sd60439, 32'sd627436, 32'sd246007, 32'sd422, 32'sd4025, 32'sd393825, 32'sd246825,
32'sd1098226, 32'sd32064, 32'sd242600, 32'sd15514, 32'sd24036, 32'sd536778, 32'sd165274, 32'sd574305, 32'sd270688, 32'sd92745,
32'sd613650, 32'sd187050, 32'sd98012, 32'sd252790, 32'sd496954, 32'sd201267, 32'sd107899, 32'sd406, 32'sd102685, 32'sd463006,
32'sd354884, 32'sd444372, 32'sd174755, 32'sd881029, 32'sd165830, 32'sd259914, 32'sd426340, 32'sd5958, 32'sd432308, 32'sd247997,
32'sd1232588, 32'sd203960, 32'sd276216, 32'sd850814, 32'sd250814, 32'sd33079, 32'sd50553, 32'sd26485, 32'sd9425, 32'sd410694,
32'sd85682, 32'sd113263, 32'sd136277, 32'sd353531, 32'sd456142, 32'sd204429, 32'sd29569, 32'sd177874, 32'sd871060, 32'sd140585,
32'sd508302, 32'sd405889, 32'sd822378, 32'sd199393, 32'sd46235, 32'sd536433, 32'sd249058, 32'sd154003, 32'sd310329, 32'sd118433,
32'sd343029, 32'sd442240, 32'sd293585, 32'sd330018, 32'sd17736, 32'sd78445, 32'sd85840, 32'sd405732, 32'sd208320, 32'sd99563,
32'sd11908, 32'sd194542, 32'sd296699, 32'sd37240, 32'sd259715, 32'sd376672, 32'sd318173, 32'sd1054545, 32'sd683856, 32'sd112668,
32'sd565731, 32'sd466743, 32'sd515420, 32'sd111224, 32'sd733842, 32'sd93165, 32'sd29607, 32'sd115400, 32'sd183750, 32'sd305216,
32'sd324283, 32'sd914172, 32'sd79242, 32'sd266962, 32'sd556846, 32'sd229122, 32'sd145543, 32'sd622810, 32'sd1315955, 32'sd212524,
32'sd307846, 32'sd720034, 32'sd9210, 32'sd33125, 32'sd384786, 32'sd283493, 32'sd19476, 32'sd406112, 32'sd378387, 32'sd351195,
32'sd288155, 32'sd115197, 32'sd125388, 32'sd403266, 32'sd271925, 32'sd695067, 32'sd131662, 32'sd106366, 32'sd62630, 32'sd230194,
32'sd34644, 32'sd629934, 32'sd25153, 32'sd587811, 32'sd612147, 32'sd260557, 32'sd32093, 32'sd694722, 32'sd159825, 32'sd186267,
32'sd388631, 32'sd386289, 32'sd165638, 32'sd448437, 32'sd18554, 32'sd215662, 32'sd324934, 32'sd395681, 32'sd10835, 32'sd304355,
32'sd49769, 32'sd584155, 32'sd678215, 32'sd63261, 32'sd116898, 32'sd402797, 32'sd351747, 32'sd81028, 32'sd61617, 32'sd32835,
32'sd229365, 32'sd305051, 32'sd481409, 32'sd330978, 32'sd333360, 32'sd35325, 32'sd923214, 32'sd49416, 32'sd177015, 32'sd312336,
32'sd39807, 32'sd546851, 32'sd677003, 32'sd242667, 32'sd5266, 32'sd15496, 32'sd704899, 32'sd917618, 32'sd182063, 32'sd467455,
32'sd76859, 32'sd543573, 32'sd589447, 32'sd36706, 32'sd2565, 32'sd83745, 32'sd61302, 32'sd288939, 32'sd117907, 32'sd217585,
32'sd202961, 32'sd468938, 32'sd80475, 32'sd558777, 32'sd231210, 32'sd37145, 32'sd1230049, 32'sd113058, 32'sd31462, 32'sd432085,
32'sd656919, 32'sd394514, 32'sd65021, 32'sd195129, 32'sd67412, 32'sd213099, 32'sd362130, 32'sd200463, 32'sd75936, 32'sd542868,
32'sd427463, 32'sd521180, 32'sd22053, 32'sd973240, 32'sd831, 32'sd524398, 32'sd744966, 32'sd805730, 32'sd725641, 32'sd1007447,
32'sd209006, 32'sd648240, 32'sd5395, 32'sd196919, 32'sd69985, 32'sd82400, 32'sd194890, 32'sd119308, 32'sd229705, 32'sd199715,
32'sd190452, 32'sd122475, 32'sd50409, 32'sd18818, 32'sd856767, 32'sd229050, 32'sd478614, 32'sd589530, 32'sd149316, 32'sd228952,
32'sd203895, 32'sd529204, 32'sd476133, 32'sd185743, 32'sd41415, 32'sd203070, 32'sd186771, 32'sd634286, 32'sd305610, 32'sd103212,
32'sd143208, 32'sd367731, 32'sd201845, 32'sd103894, 32'sd436411, 32'sd76659, 32'sd1020946, 32'sd355303, 32'sd37738, 32'sd289536,
32'sd378723, 32'sd212864, 32'sd166476, 32'sd426967, 32'sd302507, 32'sd243968, 32'sd720776, 32'sd35298, 32'sd522114, 32'sd53368,
32'sd185661, 32'sd241937, 32'sd21825, 32'sd76386, 32'sd305543, 32'sd131970, 32'sd22792, 32'sd124674, 32'sd420340, 32'sd26862,
32'sd136513, 32'sd329832, 32'sd134711, 32'sd627261, 32'sd771986, 32'sd28522, 32'sd202584, 32'sd192401, 32'sd225149, 32'sd617898,
32'sd85294, 32'sd76330, 32'sd185865, 32'sd197746, 32'sd60430, 32'sd285352, 32'sd242577, 32'sd326756, 32'sd223547, 32'sd323335,
32'sd344422, 32'sd260964, 32'sd233757, 32'sd150159, 32'sd426649, 32'sd414482, 32'sd819506, 32'sd752117, 32'sd74383, 32'sd69548,
32'sd140074, 32'sd391812, 32'sd114980, 32'sd53973, 32'sd15029, 32'sd232957, 32'sd588922, 32'sd122551, 32'sd252166, 32'sd179385,
32'sd155286, 32'sd218115, 32'sd66909, 32'sd273106, 32'sd260146, 32'sd79135, 32'sd246496, 32'sd527442, 32'sd95810, 32'sd82032,
32'sd91910, 32'sd47110, 32'sd298344, 32'sd348774, 32'sd140142, 32'sd86213, 32'sd22257, 32'sd235595, 32'sd230458, 32'sd342322,
32'sd20180, 32'sd161032, 32'sd916, 32'sd870740, 32'sd235134, 32'sd184380, 32'sd41404, 32'sd75132, 32'sd281395, 32'sd232731,
32'sd402021, 32'sd62568, 32'sd12993, 32'sd108473, 32'sd247844, 32'sd140581, 32'sd293940, 32'sd289736, 32'sd256951, 32'sd112350,
32'sd43181, 32'sd154528, 32'sd158547, 32'sd258249, 32'sd82867, 32'sd84764, 32'sd161507, 32'sd454902, 32'sd317663, 32'sd234877,
32'sd136818, 32'sd527747, 32'sd196014, 32'sd66851, 32'sd707202, 32'sd416897, 32'sd494879, 32'sd228541, 32'sd56620, 32'sd6240,
32'sd418615, 32'sd91138, 32'sd1029540, 32'sd116650, 32'sd391021, 32'sd514310, 32'sd40256, 32'sd474953, 32'sd663335, 32'sd429975,
32'sd629615, 32'sd116980, 32'sd290997, 32'sd247617, 32'sd677557, 32'sd221901, 32'sd559028, 32'sd316072, 32'sd229173, 32'sd181539,
32'sd56746, 32'sd20640, 32'sd521001, 32'sd158725, 32'sd139130, 32'sd1399986, 32'sd463396, 32'sd103308, 32'sd204926, 32'sd648079,
32'sd117343, 32'sd225653, 32'sd2431, 32'sd490370, 32'sd699331, 32'sd121727, 32'sd373, 32'sd518379, 32'sd124878, 32'sd709089,
32'sd460730, 32'sd470582, 32'sd56534, 32'sd201709, 32'sd110367, 32'sd709378, 32'sd157084, 32'sd91884, 32'sd96695, 32'sd87184,
32'sd20352, 32'sd451270, 32'sd671507, 32'sd335299, 32'sd129090, 32'sd288811, 32'sd360290, 32'sd46464, 32'sd813804, 32'sd183678,
32'sd120973, 32'sd75516, 32'sd943932, 32'sd258280, 32'sd253311, 32'sd623745, 32'sd114161, 32'sd183022, 32'sd175480, 32'sd292248,
32'sd191729, 32'sd206228, 32'sd33100, 32'sd486499, 32'sd375429, 32'sd40661, 32'sd367756, 32'sd380685, 32'sd663319, 32'sd685857,
32'sd114323, 32'sd641325, 32'sd426929, 32'sd140349, 32'sd320296, 32'sd170683, 32'sd326988, 32'sd199856, 32'sd582602, 32'sd545384,
32'sd69355, 32'sd206706, 32'sd102164, 32'sd716417, 32'sd201048, 32'sd130398, 32'sd173575, 32'sd29951, 32'sd26924, 32'sd80609,
32'sd139004, 32'sd1229692, 32'sd206382, 32'sd150398, 32'sd11782, 32'sd238667, 32'sd519714, 32'sd71238, 32'sd213619, 32'sd68543,
32'sd532266, 32'sd151877, 32'sd113360, 32'sd172094, 32'sd27078, 32'sd59509, 32'sd377424, 32'sd94758, 32'sd194888, 32'sd596676,
32'sd9564, 32'sd110535, 32'sd155265, 32'sd64270, 32'sd309666, 32'sd340589, 32'sd164281, 32'sd98389, 32'sd531933, 32'sd51557,
32'sd414158, 32'sd95796, 32'sd115734, 32'sd10822, 32'sd128803, 32'sd652453, 32'sd427475, 32'sd221201, 32'sd220732, 32'sd361136,
32'sd103898, 32'sd828737, 32'sd478968, 32'sd214239, 32'sd246829, 32'sd143090, 32'sd235045, 32'sd210168, 32'sd527934, 32'sd47057,
32'sd165694, 32'sd29855, 32'sd43602, 32'sd407278, 32'sd70273, 32'sd123747, 32'sd21586, 32'sd13106, 32'sd1095614, 32'sd631900,
32'sd199877, 32'sd561248, 32'sd74674, 32'sd268574, 32'sd318729, 32'sd1024668, 32'sd812326, 32'sd17680, 32'sd348150, 32'sd736593,
32'sd49277, 32'sd28402, 32'sd534268, 32'sd17582, 32'sd467101, 32'sd334884, 32'sd75855, 32'sd280563, 32'sd310638, 32'sd83412,
32'sd306186, 32'sd99913, 32'sd545308, 32'sd262624, 32'sd128618, 32'sd704012, 32'sd679620, 32'sd637811, 32'sd281959, 32'sd470837,
32'sd43472, 32'sd177272, 32'sd302426, 32'sd25950, 32'sd477487, 32'sd24722, 32'sd32820, 32'sd132543, 32'sd386603, 32'sd215654,
32'sd239140, 32'sd137851, 32'sd596221, 32'sd51822, 32'sd29791, 32'sd11654, 32'sd294553, 32'sd72980, 32'sd192517, 32'sd148254,
32'sd45654, 32'sd692163, 32'sd617539, 32'sd427219, 32'sd285409, 32'sd619379, 32'sd223111, 32'sd409293, 32'sd70354, 32'sd401108,
32'sd147436, 32'sd191997, 32'sd27454, 32'sd335366, 32'sd771459, 32'sd16589, 32'sd41037, 32'sd118678, 32'sd51820, 32'sd307457,
32'sd728825, 32'sd841467, 32'sd141060, 32'sd194740, 32'sd350548, 32'sd28022, 32'sd173888, 32'sd270166, 32'sd171420, 32'sd15109,
32'sd731859, 32'sd15210, 32'sd31465, 32'sd624673, 32'sd318498, 32'sd486198, 32'sd80856, 32'sd638710, 32'sd592780, 32'sd219596,
32'sd231556, 32'sd237547, 32'sd733699, 32'sd387273, 32'sd528855, 32'sd608732, 32'sd2643, 32'sd273457, 32'sd130040, 32'sd244025,
32'sd9935, 32'sd898524, 32'sd172795, 32'sd238422, 32'sd7645, 32'sd188660, 32'sd45393, 32'sd891948, 32'sd161396, 32'sd167432,
32'sd128218, 32'sd122915, 32'sd307458, 32'sd325698, 32'sd218925, 32'sd337456, 32'sd831102, 32'sd268421, 32'sd99452, 32'sd439551,
32'sd260901, 32'sd162780, 32'sd69362, 32'sd67418, 32'sd157530, 32'sd602989, 32'sd52683, 32'sd405658, 32'sd420197, 32'sd199035,
32'sd203923, 32'sd131310, 32'sd2910, 32'sd682165, 32'sd241646, 32'sd225619, 32'sd418201, 32'sd585392, 32'sd130233, 32'sd169695,
32'sd215308, 32'sd365296, 32'sd44420, 32'sd170155, 32'sd214525, 32'sd100629, 32'sd214956, 32'sd165313, 32'sd461458, 32'sd323301,
32'sd44096, 32'sd395366, 32'sd421640, 32'sd654152, 32'sd50294, 32'sd49951, 32'sd57592, 32'sd514942, 32'sd11746, 32'sd536903,
32'sd420150, 32'sd17996, 32'sd769827, 32'sd11765, 32'sd166488, 32'sd97535, 32'sd64363, 32'sd416951, 32'sd88555, 32'sd30213,
32'sd296818, 32'sd66348, 32'sd199720, 32'sd450000, 32'sd233406, 32'sd199962, 32'sd436398, 32'sd7156, 32'sd18502, 32'sd200039,
32'sd341707, 32'sd95935, 32'sd208161, 32'sd145785, 32'sd1408942, 32'sd375521, 32'sd50977, 32'sd641982, 32'sd249066, 32'sd312543,
32'sd471541, 32'sd51586, 32'sd652135, 32'sd145717, 32'sd32414, 32'sd233094, 32'sd470012, 32'sd501510, 32'sd884194, 32'sd1110,
32'sd95476, 32'sd4197, 32'sd431144, 32'sd297479, 32'sd449974, 32'sd53841, 32'sd152627, 32'sd422667, 32'sd464403, 32'sd100024,
32'sd408777, 32'sd218623, 32'sd212111, 32'sd415728, 32'sd242717, 32'sd6169, 32'sd5217, 32'sd193475, 32'sd414837, 32'sd308738,
32'sd13007, 32'sd504894, 32'sd283109, 32'sd177739, 32'sd246880, 32'sd16649, 32'sd229145, 32'sd42447, 32'sd133785, 32'sd494596,
32'sd670614, 32'sd5267, 32'sd252097, 32'sd786473, 32'sd224342, 32'sd147187, 32'sd32232, 32'sd43409, 32'sd401257, 32'sd891121,
32'sd266669, 32'sd64797, 32'sd76857, 32'sd157124, 32'sd27060, 32'sd148875, 32'sd160478, 32'sd27393, 32'sd91457, 32'sd203543,
32'sd532612, 32'sd84245, 32'sd105832, 32'sd19317, 32'sd332501, 32'sd142817, 32'sd586571, 32'sd276767, 32'sd87098, 32'sd354535,
32'sd48142, 32'sd143179, 32'sd31458, 32'sd174165, 32'sd746663, 32'sd62393, 32'sd288726, 32'sd831300, 32'sd24328, 32'sd445776,
32'sd172324, 32'sd532552, 32'sd245070, 32'sd6325, 32'sd164324, 32'sd81300, 32'sd145792, 32'sd777610, 32'sd210058, 32'sd31215,
32'sd267995, 32'sd199945, 32'sd446714, 32'sd625128, 32'sd15325, 32'sd95482, 32'sd198014, 32'sd146684, 32'sd111954, 32'sd604040,
32'sd99053, 32'sd306519, 32'sd123660, 32'sd74408, 32'sd107382, 32'sd385489, 32'sd99915, 32'sd491178, 32'sd319144, 32'sd9551,
32'sd198641, 32'sd109386, 32'sd47144, 32'sd23508, 32'sd127148, 32'sd901162, 32'sd20364, 32'sd513387, 32'sd421989, 32'sd219200,
32'sd297273, 32'sd302776, 32'sd16488, 32'sd77034, 32'sd114753, 32'sd236392, 32'sd74885, 32'sd247120, 32'sd859131, 32'sd219901,
32'sd134252, 32'sd141072, 32'sd173047, 32'sd406691, 32'sd159883, 32'sd35789, 32'sd275442, 32'sd449080, 32'sd99837, 32'sd518683,
32'sd560752, 32'sd464838, 32'sd159437, 32'sd287213, 32'sd35404, 32'sd10668, 32'sd131879, 32'sd79058, 32'sd671627, 32'sd740649,
32'sd680074, 32'sd492157, 32'sd240219, 32'sd93105, 32'sd576388, 32'sd40357, 32'sd216732, 32'sd57402, 32'sd127205, 32'sd423699,
32'sd213562, 32'sd304474, 32'sd9795, 32'sd24031, 32'sd763906, 32'sd84640, 32'sd369806, 32'sd355565, 32'sd473155, 32'sd137086,
32'sd79813, 32'sd213826, 32'sd74678, 32'sd400836, 32'sd68919, 32'sd247206, 32'sd229131, 32'sd261692, 32'sd977344, 32'sd11842,
32'sd249908, 32'sd243220, 32'sd98654, 32'sd682315, 32'sd351500, 32'sd331011, 32'sd134664, 32'sd67833, 32'sd1386263, 32'sd166867,
32'sd511515, 32'sd175029, 32'sd332066, 32'sd143061, 32'sd62249, 32'sd61753, 32'sd76080, 32'sd140176, 32'sd205, 32'sd393118,
32'sd555280, 32'sd308740, 32'sd719456, 32'sd435632, 32'sd521271, 32'sd19288, 32'sd109595, 32'sd128102, 32'sd245895, 32'sd1084422,
32'sd651304, 32'sd511831, 32'sd543680, 32'sd469406, 32'sd767472, 32'sd1179057, 32'sd923320, 32'sd82586, 32'sd519257, 32'sd1045080,
32'sd649676, 32'sd36061, 32'sd458970, 32'sd42921, 32'sd188437, 32'sd124359, 32'sd218569, 32'sd464386, 32'sd80368, 32'sd161068,
32'sd33381, 32'sd498654, 32'sd409659, 32'sd476054, 32'sd327157, 32'sd483692, 32'sd259550, 32'sd321357, 32'sd110188, 32'sd28080,
32'sd280151, 32'sd513088, 32'sd315782, 32'sd379012, 32'sd438783, 32'sd24113, 32'sd12308, 32'sd79713, 32'sd271324, 32'sd48180,
32'sd210320, 32'sd45821, 32'sd437106, 32'sd664627, 32'sd54384, 32'sd62077, 32'sd111864, 32'sd239809, 32'sd447989, 32'sd355085,
32'sd854937, 32'sd321412, 32'sd53603, 32'sd224618, 32'sd101915, 32'sd319059, 32'sd633700, 32'sd269992, 32'sd411988, 32'sd304384,
32'sd288612, 32'sd288267, 32'sd368512, 32'sd119419, 32'sd728783, 32'sd43821, 32'sd1274471, 32'sd273210, 32'sd241598, 32'sd110591,
32'sd17197, 32'sd550200, 32'sd317574, 32'sd126652, 32'sd220453, 32'sd16657, 32'sd475978, 32'sd246214, 32'sd127105, 32'sd17142,
32'sd138138, 32'sd214950, 32'sd590062, 32'sd83130, 32'sd15347, 32'sd120159, 32'sd432561, 32'sd953968, 32'sd496585, 32'sd150670,
32'sd761374, 32'sd340337, 32'sd800886, 32'sd223510, 32'sd538991, 32'sd84034, 32'sd626878, 32'sd213007, 32'sd73086, 32'sd471021,
32'sd4617, 32'sd164226, 32'sd813041, 32'sd401915, 32'sd388370, 32'sd52302, 32'sd325095, 32'sd61411, 32'sd322429, 32'sd511653,
32'sd19031, 32'sd78102, 32'sd978760, 32'sd33964, 32'sd115945, 32'sd14652, 32'sd530746, 32'sd31023, 32'sd106724, 32'sd299825,
32'sd45604, 32'sd24759, 32'sd84274, 32'sd695437, 32'sd144603, 32'sd289503, 32'sd539859, 32'sd877412, 32'sd373612, 32'sd244606,
32'sd136110, 32'sd650907, 32'sd680841, 32'sd198497, 32'sd451515, 32'sd237169, 32'sd646228, 32'sd291120, 32'sd229204, 32'sd57090,
32'sd194969, 32'sd159236, 32'sd188569, 32'sd1035670, 32'sd16856, 32'sd74004, 32'sd476629, 32'sd393013, 32'sd38608, 32'sd285153,
32'sd207867, 32'sd5458, 32'sd330237, 32'sd97300, 32'sd1090740, 32'sd10648, 32'sd325934, 32'sd322136, 32'sd291930, 32'sd778482,
32'sd714714, 32'sd308493, 32'sd83916, 32'sd257364, 32'sd291186, 32'sd702714, 32'sd245135, 32'sd608492, 32'sd483380, 32'sd743620,
32'sd1106434, 32'sd3051, 32'sd246316, 32'sd309983, 32'sd389824, 32'sd759137, 32'sd136489, 32'sd343531, 32'sd37407, 32'sd140031,
32'sd400932, 32'sd581731, 32'sd204190, 32'sd320424, 32'sd564318, 32'sd239979, 32'sd172305, 32'sd486850, 32'sd295339, 32'sd608834,
32'sd359984, 32'sd12624, 32'sd92214, 32'sd43710, 32'sd102057, 32'sd148244, 32'sd63396, 32'sd295116, 32'sd287337, 32'sd111078,
32'sd32531, 32'sd828054, 32'sd405104, 32'sd308875, 32'sd78957, 32'sd271647, 32'sd680927, 32'sd906466, 32'sd217958, 32'sd22551,
32'sd144226, 32'sd130143, 32'sd165872, 32'sd147584, 32'sd878094, 32'sd582842, 32'sd273394, 32'sd752162, 32'sd12740, 32'sd411686,
32'sd427851, 32'sd298072, 32'sd77324, 32'sd367067, 32'sd620040, 32'sd255493, 32'sd47904, 32'sd175820, 32'sd80052, 32'sd50656,
32'sd278998, 32'sd58102, 32'sd160987, 32'sd293157, 32'sd471579, 32'sd715364, 32'sd173197, 32'sd19644, 32'sd334796, 32'sd281064,
32'sd206950, 32'sd29229, 32'sd330232, 32'sd222279, 32'sd655184, 32'sd338005, 32'sd394818, 32'sd470307, 32'sd145780, 32'sd707989,
32'sd563949, 32'sd580714, 32'sd1007745, 32'sd28844, 32'sd811342, 32'sd183672, 32'sd35057, 32'sd846631, 32'sd235978, 32'sd8698,
32'sd998163, 32'sd681919, 32'sd46915, 32'sd492047, 32'sd272831, 32'sd230090, 32'sd125399, 32'sd854041, 32'sd337295, 32'sd204334,
32'sd389491, 32'sd33614, 32'sd491091, 32'sd689251, 32'sd234540, 32'sd118759, 32'sd858402, 32'sd113995, 32'sd331, 32'sd56628,
32'sd252011, 32'sd152667, 32'sd263310, 32'sd57045, 32'sd224235, 32'sd230100, 32'sd14428, 32'sd16488, 32'sd417308, 32'sd66234,
32'sd1435, 32'sd8417, 32'sd10291, 32'sd443479, 32'sd152798, 32'sd682131, 32'sd234360, 32'sd84954, 32'sd164413, 32'sd84904,
32'sd96561, 32'sd434212, 32'sd76130, 32'sd241068, 32'sd213820, 32'sd469442, 32'sd355930, 32'sd13338, 32'sd552037, 32'sd119543,
32'sd65808, 32'sd452553, 32'sd76265, 32'sd559184, 32'sd196387, 32'sd254539, 32'sd3928, 32'sd206634, 32'sd152030, 32'sd48111,
32'sd67155, 32'sd584579, 32'sd23770, 32'sd312556, 32'sd367654, 32'sd638744, 32'sd610015, 32'sd84237, 32'sd8406, 32'sd250156,
32'sd226600, 32'sd372604, 32'sd289740, 32'sd250794, 32'sd46362, 32'sd48836, 32'sd558916, 32'sd494999, 32'sd388036, 32'sd479246,
32'sd700276, 32'sd157197, 32'sd268311, 32'sd482940, 32'sd184126, 32'sd300668, 32'sd114352, 32'sd262718, 32'sd19197, 32'sd982670,
32'sd199371, 32'sd1006042, 32'sd314887, 32'sd210470, 32'sd356250, 32'sd170663, 32'sd19393, 32'sd106020, 32'sd55600, 32'sd256550,
32'sd33925, 32'sd94411, 32'sd482248, 32'sd146262, 32'sd479932, 32'sd122069, 32'sd16893, 32'sd199023, 32'sd620581, 32'sd128783,
32'sd257930, 32'sd99448, 32'sd321556, 32'sd157634, 32'sd449507, 32'sd259299, 32'sd235566, 32'sd69741, 32'sd853102, 32'sd571224,
32'sd352314, 32'sd517171, 32'sd9563, 32'sd462980, 32'sd516204, 32'sd40467, 32'sd68603, 32'sd243740, 32'sd167870, 32'sd145392,
32'sd281907, 32'sd578475, 32'sd44657, 32'sd155977, 32'sd386218, 32'sd590818, 32'sd46920, 32'sd178433, 32'sd152837, 32'sd164004,
32'sd765624, 32'sd23683, 32'sd935802, 32'sd1501257, 32'sd27924, 32'sd530411, 32'sd42879, 32'sd485562, 32'sd265172, 32'sd217041,
32'sd769067, 32'sd76159, 32'sd397106, 32'sd495807, 32'sd92154, 32'sd169065, 32'sd630551, 32'sd368382, 32'sd1193830, 32'sd273702,
32'sd117934, 32'sd50485, 32'sd467606, 32'sd632001, 32'sd24334, 32'sd207166, 32'sd647954, 32'sd6702, 32'sd10767, 32'sd3601,
32'sd120023, 32'sd246331, 32'sd312524, 32'sd62007, 32'sd669854, 32'sd100973, 32'sd525400, 32'sd99254, 32'sd131760, 32'sd329722,
32'sd171640, 32'sd236333, 32'sd214615, 32'sd552744, 32'sd5878, 32'sd214014, 32'sd510854, 32'sd16076, 32'sd157289, 32'sd188740,
32'sd345307, 32'sd56151, 32'sd112670, 32'sd235635, 32'sd355302, 32'sd276030, 32'sd86261, 32'sd156358, 32'sd51747, 32'sd178153,
32'sd106176, 32'sd274494, 32'sd677756, 32'sd805211, 32'sd48498, 32'sd178903, 32'sd626822, 32'sd264340, 32'sd429378, 32'sd346515,
32'sd63053, 32'sd310301, 32'sd476356, 32'sd58393, 32'sd104704, 32'sd240321, 32'sd32071, 32'sd50361, 32'sd266150, 32'sd901935,
32'sd151584, 32'sd484864, 32'sd88306, 32'sd43374, 32'sd226343, 32'sd339597, 32'sd826500, 32'sd386765, 32'sd469216, 32'sd22886,
32'sd73721, 32'sd69386, 32'sd213851, 32'sd81967, 32'sd276499, 32'sd507264, 32'sd262817, 32'sd28249, 32'sd518035, 32'sd139621,
32'sd36265, 32'sd58769, 32'sd259635, 32'sd507616, 32'sd242375, 32'sd366683, 32'sd181549, 32'sd6045, 32'sd2495, 32'sd602589,
32'sd740501, 32'sd332631, 32'sd16726, 32'sd803799, 32'sd323135, 32'sd57693, 32'sd188276, 32'sd1094485, 32'sd222851, 32'sd632820,
32'sd310687, 32'sd169872, 32'sd338291, 32'sd42380, 32'sd127832, 32'sd252602, 32'sd493331, 32'sd591223, 32'sd231786, 32'sd237147,
32'sd170551, 32'sd10957, 32'sd110948, 32'sd222540, 32'sd789708, 32'sd86427, 32'sd888714, 32'sd325812, 32'sd359538, 32'sd619385,
32'sd84054, 32'sd399992, 32'sd174672, 32'sd743786, 32'sd73369, 32'sd912820, 32'sd51555, 32'sd333060, 32'sd110750, 32'sd150803,
32'sd242049, 32'sd654153, 32'sd135887, 32'sd66849, 32'sd184090, 32'sd198564, 32'sd415591, 32'sd385350, 32'sd234595, 32'sd68672,
32'sd351987, 32'sd281648, 32'sd395505, 32'sd277753, 32'sd155820, 32'sd100018, 32'sd125988, 32'sd115397, 32'sd477582, 32'sd142937,
32'sd260221, 32'sd63813, 32'sd783735, 32'sd518496, 32'sd5454, 32'sd723211, 32'sd86373, 32'sd13494, 32'sd71514, 32'sd181488,
32'sd575292, 32'sd72725, 32'sd302225, 32'sd116727, 32'sd26203, 32'sd31058, 32'sd284628, 32'sd532268, 32'sd197669, 32'sd205634,
32'sd59890, 32'sd143481, 32'sd168568, 32'sd180464, 32'sd231822, 32'sd110292, 32'sd48534, 32'sd191198, 32'sd409583, 32'sd83186,
32'sd513824, 32'sd172870, 32'sd9125, 32'sd857251, 32'sd842159, 32'sd107385, 32'sd1012409, 32'sd515287, 32'sd304167, 32'sd54451,
32'sd535005, 32'sd540264, 32'sd75764, 32'sd23046, 32'sd516876, 32'sd12488, 32'sd54662, 32'sd161558, 32'sd641253, 32'sd667052,
32'sd176104, 32'sd789680, 32'sd131427, 32'sd14741, 32'sd327531, 32'sd346070, 32'sd613129, 32'sd82120, 32'sd28887, 32'sd388538,
32'sd235772, 32'sd418454, 32'sd54040, 32'sd49028, 32'sd173430, 32'sd797602, 32'sd593370, 32'sd632267, 32'sd457020, 32'sd905307,
32'sd536938, 32'sd6787, 32'sd103193, 32'sd38239, 32'sd226114, 32'sd73200, 32'sd22916, 32'sd178913, 32'sd51618, 32'sd410479,
32'sd191600, 32'sd1059770, 32'sd7034, 32'sd325647, 32'sd50306, 32'sd131233, 32'sd297092, 32'sd363478, 32'sd176699, 32'sd110752,
32'sd3758, 32'sd153012, 32'sd333672, 32'sd363032, 32'sd652261, 32'sd492742, 32'sd410426, 32'sd360091, 32'sd780990, 32'sd338198,
32'sd134544, 32'sd550335, 32'sd201876, 32'sd435096, 32'sd149966, 32'sd284739, 32'sd624345, 32'sd466547, 32'sd417448, 32'sd314481,
32'sd106251, 32'sd94513, 32'sd85832, 32'sd348168, 32'sd587856, 32'sd5105, 32'sd212234, 32'sd372644, 32'sd15021, 32'sd175211,
32'sd7467, 32'sd84840, 32'sd516229, 32'sd245930, 32'sd88200, 32'sd332046, 32'sd19544, 32'sd161622, 32'sd598514, 32'sd111289,
32'sd375036, 32'sd603279, 32'sd216991, 32'sd262114, 32'sd656020, 32'sd458393, 32'sd20012, 32'sd802657, 32'sd190659, 32'sd274343,
32'sd62157, 32'sd414241, 32'sd361871, 32'sd258270, 32'sd251997, 32'sd225609, 32'sd397454, 32'sd395666, 32'sd373374, 32'sd55013,
32'sd311677, 32'sd1700, 32'sd222468, 32'sd592648, 32'sd310903, 32'sd147901, 32'sd247078, 32'sd26887, 32'sd596084, 32'sd198256,
32'sd227344, 32'sd698990, 32'sd360378, 32'sd141354, 32'sd172915, 32'sd220048, 32'sd67760, 32'sd143512, 32'sd380035, 32'sd229979,
32'sd424654, 32'sd1413509, 32'sd94367, 32'sd272802, 32'sd928591, 32'sd314039, 32'sd748576, 32'sd270782, 32'sd95370, 32'sd184737,
32'sd127589, 32'sd151073, 32'sd1031407, 32'sd349687, 32'sd15012, 32'sd371290, 32'sd172301, 32'sd32295, 32'sd197257, 32'sd95030,
32'sd313427, 32'sd187341, 32'sd251816, 32'sd812866, 32'sd159421, 32'sd69351, 32'sd327137, 32'sd161051, 32'sd292007, 32'sd59963,
32'sd147370, 32'sd434580, 32'sd61783, 32'sd41147, 32'sd561905, 32'sd339374, 32'sd106268, 32'sd636902, 32'sd712106, 32'sd429455,
32'sd854630, 32'sd305739, 32'sd190679, 32'sd676579, 32'sd477620, 32'sd793, 32'sd83565, 32'sd402713, 32'sd73640, 32'sd237465,
32'sd25214, 32'sd185231, 32'sd5884, 32'sd203736, 32'sd77196, 32'sd722022, 32'sd148562, 32'sd386915, 32'sd648809, 32'sd114291,
32'sd162359, 32'sd282479, 32'sd25942, 32'sd72044, 32'sd59712, 32'sd806511, 32'sd152260, 32'sd65725, 32'sd439834, 32'sd80002,
32'sd289092, 32'sd67186, 32'sd1213741, 32'sd105156, 32'sd107315, 32'sd295819, 32'sd303355, 32'sd288619, 32'sd211772, 32'sd240984,
32'sd507682, 32'sd295766, 32'sd463502, 32'sd333906, 32'sd6595, 32'sd1077866, 32'sd196108, 32'sd341805, 32'sd157718, 32'sd371983,
32'sd641555, 32'sd69860, 32'sd348582, 32'sd103193, 32'sd734645, 32'sd334642, 32'sd626613, 32'sd175179, 32'sd1038207, 32'sd1172753,
32'sd312768, 32'sd97599, 32'sd787500, 32'sd663554, 32'sd724547, 32'sd132823, 32'sd509329, 32'sd74613, 32'sd116149, 32'sd145359,
32'sd458773, 32'sd368568, 32'sd194309, 32'sd130566, 32'sd684820, 32'sd11923, 32'sd65160, 32'sd906766, 32'sd191406, 32'sd521927,
32'sd194221, 32'sd313992, 32'sd53165, 32'sd239091, 32'sd227575, 32'sd32565, 32'sd329521, 32'sd110011, 32'sd40101, 32'sd556150,
32'sd85397, 32'sd101978, 32'sd251234, 32'sd9150, 32'sd460604, 32'sd500159, 32'sd248460, 32'sd2023, 32'sd622389, 32'sd235159,
32'sd267713, 32'sd71018, 32'sd65895, 32'sd265179, 32'sd33994, 32'sd40968, 32'sd117659, 32'sd425634, 32'sd73499, 32'sd20342,
32'sd126277, 32'sd202547, 32'sd31884, 32'sd785578, 32'sd82752, 32'sd332038, 32'sd743285, 32'sd8571, 32'sd517190, 32'sd535553,
32'sd880979, 32'sd13917, 32'sd212758, 32'sd32120, 32'sd25395, 32'sd275869, 32'sd17875, 32'sd84005, 32'sd69122, 32'sd312128,
32'sd541034, 32'sd589209, 32'sd184562, 32'sd612432, 32'sd317490, 32'sd217969, 32'sd26601, 32'sd68543, 32'sd17328, 32'sd42571,
32'sd472344, 32'sd1229, 32'sd212567, 32'sd425214, 32'sd39842, 32'sd75379, 32'sd1179149, 32'sd641920, 32'sd240620, 32'sd401026,
32'sd449792, 32'sd177939, 32'sd302111, 32'sd20831, 32'sd234065, 32'sd2392, 32'sd220851, 32'sd271356, 32'sd73312, 32'sd359240,
32'sd307260, 32'sd727446, 32'sd396729, 32'sd156195, 32'sd65725, 32'sd492573, 32'sd145945, 32'sd122237, 32'sd325466, 32'sd94567,
32'sd631069, 32'sd27775, 32'sd350874, 32'sd138175, 32'sd398772, 32'sd107934, 32'sd7594, 32'sd89330, 32'sd143880, 32'sd520807,
32'sd45456, 32'sd386961, 32'sd70368, 32'sd83031, 32'sd1133695, 32'sd296903, 32'sd224660, 32'sd421607, 32'sd22567, 32'sd91637,
32'sd169710, 32'sd714665, 32'sd666720, 32'sd16322, 32'sd391230, 32'sd210636, 32'sd29629, 32'sd32949, 32'sd14561, 32'sd38799,
32'sd484613, 32'sd435020, 32'sd1006351, 32'sd94682, 32'sd6815, 32'sd29878, 32'sd28692, 32'sd251977, 32'sd212476, 32'sd540402,
32'sd94662, 32'sd39291, 32'sd597660, 32'sd45983, 32'sd260923, 32'sd460228, 32'sd8418, 32'sd128100, 32'sd613921, 32'sd417443,
32'sd387009, 32'sd125877, 32'sd194295, 32'sd22016, 32'sd204017, 32'sd80075, 32'sd65449, 32'sd541721, 32'sd128873, 32'sd227953,
32'sd71707, 32'sd170430, 32'sd306280, 32'sd79116, 32'sd245812, 32'sd131611, 32'sd108758, 32'sd386761, 32'sd803413, 32'sd204806,
32'sd54471, 32'sd452218, 32'sd22178, 32'sd376254, 32'sd1003991, 32'sd236688, 32'sd43320, 32'sd228556, 32'sd269647, 32'sd147007,
32'sd830695, 32'sd418924, 32'sd539283, 32'sd30482, 32'sd844646, 32'sd539074, 32'sd111008, 32'sd88007, 32'sd75231, 32'sd395298,
32'sd301752, 32'sd669483, 32'sd302034, 32'sd448233, 32'sd47002, 32'sd579543, 32'sd610178, 32'sd39244, 32'sd238832, 32'sd92346,
32'sd305346, 32'sd80070, 32'sd402393, 32'sd911124, 32'sd317383, 32'sd387758, 32'sd1105881, 32'sd442436, 32'sd124442, 32'sd309553,
32'sd24195, 32'sd179709, 32'sd276291, 32'sd783, 32'sd1059901, 32'sd75130, 32'sd303409, 32'sd759470, 32'sd275090, 32'sd164352,
32'sd173528, 32'sd313198, 32'sd303976, 32'sd40944, 32'sd277814, 32'sd1075156, 32'sd128662, 32'sd36800, 32'sd68197, 32'sd670192,
32'sd134105, 32'sd969399, 32'sd308824, 32'sd384427, 32'sd6502, 32'sd385164, 32'sd255850, 32'sd26380, 32'sd174748, 32'sd434291,
32'sd26517, 32'sd1119295, 32'sd921168, 32'sd611567, 32'sd690718, 32'sd45836, 32'sd308012, 32'sd904811, 32'sd268482, 32'sd535179,
32'sd45762, 32'sd258954, 32'sd751245, 32'sd8360, 32'sd773995, 32'sd119000, 32'sd259762, 32'sd18883, 32'sd77176, 32'sd332498,
32'sd547595, 32'sd19786, 32'sd263097, 32'sd498401, 32'sd65417, 32'sd406031, 32'sd77059, 32'sd210435, 32'sd270750, 32'sd714594,
32'sd72858, 32'sd14859, 32'sd69556, 32'sd859275, 32'sd79866, 32'sd142690, 32'sd276395, 32'sd463786, 32'sd122166, 32'sd879737,
32'sd26867, 32'sd208910, 32'sd114407, 32'sd91472, 32'sd185682, 32'sd27029, 32'sd381648, 32'sd94756, 32'sd583499, 32'sd19135,
32'sd307389, 32'sd3590, 32'sd312646, 32'sd345964, 32'sd584493, 32'sd504968, 32'sd370942, 32'sd135135, 32'sd422784, 32'sd42139,
32'sd475373, 32'sd426832, 32'sd146378, 32'sd275740, 32'sd90514, 32'sd455184, 32'sd199453, 32'sd66462, 32'sd132930, 32'sd52236,
32'sd606902, 32'sd43824, 32'sd23914, 32'sd527600, 32'sd72611, 32'sd37606, 32'sd535852, 32'sd541107, 32'sd89995, 32'sd132593,
32'sd127003, 32'sd15184, 32'sd471334, 32'sd13456, 32'sd23719, 32'sd88426, 32'sd128272, 32'sd394028, 32'sd205913, 32'sd320389,
32'sd255674, 32'sd204962, 32'sd18984, 32'sd50599, 32'sd7807, 32'sd205718, 32'sd90860, 32'sd47236, 32'sd107262, 32'sd1106421,
32'sd59760, 32'sd26437, 32'sd134965, 32'sd231497, 32'sd677629, 32'sd245763, 32'sd138487, 32'sd717642, 32'sd296622, 32'sd426015,
32'sd470031, 32'sd74161, 32'sd85997, 32'sd152290, 32'sd115453, 32'sd226038, 32'sd346261, 32'sd375316, 32'sd59759, 32'sd9438,
32'sd153707, 32'sd239927, 32'sd323800, 32'sd292508, 32'sd66624, 32'sd494054, 32'sd136146, 32'sd203591, 32'sd174963, 32'sd152516,
32'sd66369, 32'sd278017, 32'sd207903, 32'sd590886, 32'sd38808, 32'sd77321, 32'sd211380, 32'sd90220, 32'sd522162, 32'sd672418,
32'sd1184111, 32'sd100306, 32'sd794, 32'sd105719, 32'sd346988, 32'sd574385, 32'sd15762, 32'sd150163, 32'sd357372, 32'sd369946,
32'sd265254, 32'sd490322, 32'sd242316, 32'sd74252, 32'sd98159, 32'sd322140, 32'sd371111, 32'sd132580, 32'sd286732, 32'sd995925,
32'sd811684, 32'sd241483, 32'sd551619, 32'sd274351, 32'sd17022, 32'sd132664, 32'sd88316, 32'sd46700, 32'sd58669, 32'sd35154,
32'sd342580, 32'sd91192, 32'sd125149, 32'sd77208, 32'sd944798, 32'sd433971, 32'sd81791, 32'sd490964, 32'sd205505, 32'sd16164,
32'sd257615, 32'sd244158, 32'sd91186, 32'sd205980, 32'sd811293, 32'sd221224, 32'sd542869, 32'sd355328, 32'sd181040, 32'sd95663,
32'sd184420, 32'sd767242, 32'sd154693, 32'sd512885, 32'sd120738, 32'sd361240, 32'sd6740, 32'sd38656, 32'sd63803, 32'sd852119,
32'sd213632, 32'sd181001

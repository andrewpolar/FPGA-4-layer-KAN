32'sd1336, 32'sd244, 32'sd1060, 32'sd922, 32'sd1770, 32'sd564,
32'sd445, 32'sd1826, 32'sd1720, 32'sd487, 32'sd1526, 32'sd121,
32'sd1366, 32'sd911, 32'sd1977, 32'sd1181, 32'sd588, 32'sd1715,
32'sd153, 32'sd1961, 32'sd1308, 32'sd714, 32'sd1710, 32'sd1154,
32'sd1499, 32'sd1229, 32'sd139, 32'sd648, 32'sd312, 32'sd1308,
32'sd665, 32'sd486, 32'sd1405, 32'sd642, 32'sd1737, 32'sd1282,
32'sd477, 32'sd845, 32'sd1349, 32'sd1155, 32'sd1430, 32'sd1821,
32'sd769, 32'sd1090, 32'sd1601, 32'sd1884, 32'sd1647, 32'sd1501,
32'sd475, 32'sd603, 32'sd1904, 32'sd907, 32'sd1006, 32'sd1945,
32'sd1367, 32'sd461, 32'sd501, 32'sd1124, 32'sd1635, 32'sd1026,
32'sd707, 32'sd1572, 32'sd658, 32'sd1434, 32'sd673, 32'sd1708,
32'sd1673, 32'sd1138, 32'sd1150, 32'sd786, 32'sd464, 32'sd1618,
32'sd1457, 32'sd1896, 32'sd1316, 32'sd1165, 32'sd1113, 32'sd1628,
32'sd1188, 32'sd1522, 32'sd123, 32'sd406, 32'sd1421, 32'sd1748,
32'sd1116, 32'sd993, 32'sd250, 32'sd1924, 32'sd125, 32'sd1049,
32'sd628, 32'sd1531, 32'sd1996, 32'sd1155, 32'sd528, 32'sd216,
32'sd299, 32'sd316, 32'sd130, 32'sd1021, 32'sd749, 32'sd993,
32'sd1636, 32'sd514, 32'sd513, 32'sd167, 32'sd1876, 32'sd792,
32'sd1979, 32'sd205, 32'sd120, 32'sd1532, 32'sd1592, 32'sd730,
32'sd1402, 32'sd1565, 32'sd1080, 32'sd1013, 32'sd611, 32'sd727,
32'sd1363, 32'sd1290, 32'sd1577, 32'sd912, 32'sd1004, 32'sd577,
32'sd1977, 32'sd357, 32'sd1043, 32'sd1546, 32'sd1376, 32'sd1844,
32'sd917, 32'sd472, 32'sd596, 32'sd1415, 32'sd1894, 32'sd1026,
32'sd1406, 32'sd129, 32'sd1354, 32'sd978, 32'sd167, 32'sd1074,
32'sd1822, 32'sd514, 32'sd896, 32'sd1360, 32'sd1004, 32'sd1225,
32'sd357, 32'sd1054, 32'sd788, 32'sd1662, 32'sd720, 32'sd500,
32'sd381, 32'sd561, 32'sd1612, 32'sd1944, 32'sd1094, 32'sd1350,
32'sd1799, 32'sd1414, 32'sd1610, 32'sd1978, 32'sd1296, 32'sd1515,
32'sd227, 32'sd1180, 32'sd1596, 32'sd1021, 32'sd820, 32'sd656,
32'sd994, 32'sd1034, 32'sd250, 32'sd1238, 32'sd391, 32'sd1840,
32'sd817, 32'sd424, 32'sd767, 32'sd881, 32'sd190, 32'sd1863,
32'sd551, 32'sd680, 32'sd473, 32'sd986, 32'sd834, 32'sd1050,
32'sd1685, 32'sd1586, 32'sd1573, 32'sd119, 32'sd1627, 32'sd1191,
32'sd464, 32'sd1588, 32'sd1352, 32'sd1886, 32'sd1119, 32'sd1491,
32'sd1004, 32'sd1933, 32'sd1330, 32'sd550, 32'sd1028, 32'sd432,
32'sd1125, 32'sd1634, 32'sd1847, 32'sd394, 32'sd966, 32'sd1617,
32'sd1310, 32'sd1935, 32'sd1246, 32'sd591, 32'sd587, 32'sd765,
32'sd1543, 32'sd897, 32'sd1128, 32'sd1371, 32'sd654, 32'sd629,
32'sd1748, 32'sd1122, 32'sd122, 32'sd264, 32'sd657, 32'sd1733,
32'sd1979, 32'sd480, 32'sd1022, 32'sd1225, 32'sd1210, 32'sd1814,
32'sd134, 32'sd805, 32'sd1793, 32'sd1873, 32'sd330, 32'sd1605,
32'sd1309, 32'sd586, 32'sd1784, 32'sd1520, 32'sd386, 32'sd900,
32'sd850, 32'sd1548, 32'sd1143, 32'sd1551, 32'sd998, 32'sd367,
32'sd1518, 32'sd1400, 32'sd1197, 32'sd182, 32'sd1124, 32'sd1038,
32'sd889, 32'sd442, 32'sd600, 32'sd184, 32'sd176, 32'sd906,
32'sd1651, 32'sd1644, 32'sd1353, 32'sd684, 32'sd561, 32'sd547,
32'sd1363, 32'sd167, 32'sd1561, 32'sd571, 32'sd1107, 32'sd1583,
32'sd1708, 32'sd1440, 32'sd720, 32'sd1211, 32'sd382, 32'sd1972,
32'sd1589, 32'sd1267, 32'sd1776, 32'sd1922, 32'sd1657, 32'sd1025,
32'sd1049, 32'sd1909, 32'sd922, 32'sd1525, 32'sd723, 32'sd976,
32'sd1108, 32'sd854, 32'sd1942, 32'sd1187, 32'sd1868, 32'sd1774,
32'sd1759, 32'sd598, 32'sd745, 32'sd1399, 32'sd1645, 32'sd1104,
32'sd822, 32'sd355, 32'sd114, 32'sd1814, 32'sd316, 32'sd1585,
32'sd1415, 32'sd921, 32'sd1508, 32'sd1060, 32'sd846, 32'sd1434,
32'sd659, 32'sd1003, 32'sd1322, 32'sd735, 32'sd1817, 32'sd1108,
32'sd1556, 32'sd254, 32'sd1992, 32'sd1490, 32'sd1967, 32'sd1773,
32'sd1763, 32'sd259, 32'sd1897, 32'sd917, 32'sd1442, 32'sd1124,
32'sd1722, 32'sd1883, 32'sd735, 32'sd1248, 32'sd1081, 32'sd256,
32'sd824, 32'sd1801, 32'sd1755, 32'sd409, 32'sd637, 32'sd644,
32'sd1999, 32'sd968, 32'sd1383, 32'sd1524, 32'sd1883, 32'sd371,
32'sd1431, 32'sd773, 32'sd1170, 32'sd872, 32'sd1276, 32'sd1505,
32'sd177, 32'sd1426, 32'sd1616, 32'sd266, 32'sd1121, 32'sd245,
32'sd700, 32'sd344, 32'sd1271, 32'sd1463, 32'sd1995, 32'sd1154,
32'sd832, 32'sd1415, 32'sd948, 32'sd106, 32'sd341, 32'sd1241,
32'sd828, 32'sd913, 32'sd1838, 32'sd124, 32'sd710, 32'sd935,
32'sd1024, 32'sd623, 32'sd458, 32'sd1077, 32'sd645, 32'sd1883,
32'sd940, 32'sd1031, 32'sd1902, 32'sd1002, 32'sd278, 32'sd534,
32'sd522, 32'sd1104, 32'sd1184, 32'sd1705, 32'sd1946, 32'sd1057,
32'sd319, 32'sd1511, 32'sd1443, 32'sd326, 32'sd1540, 32'sd143,
32'sd1069, 32'sd1074, 32'sd1504, 32'sd565, 32'sd1867, 32'sd1882,
32'sd520, 32'sd1596, 32'sd1294, 32'sd485, 32'sd1430, 32'sd1606,
32'sd882, 32'sd438, 32'sd1934, 32'sd220, 32'sd332, 32'sd985,
32'sd190, 32'sd674, 32'sd1017, 32'sd317, 32'sd531, 32'sd578,
32'sd1941, 32'sd362, 32'sd1873, 32'sd405, 32'sd141, 32'sd1018,
32'sd160, 32'sd353, 32'sd735, 32'sd741, 32'sd1489, 32'sd1925,
32'sd225, 32'sd402, 32'sd703, 32'sd1696, 32'sd467, 32'sd1075,
32'sd658, 32'sd1801, 32'sd1091, 32'sd518, 32'sd945, 32'sd1065,
32'sd125, 32'sd941, 32'sd1240, 32'sd1293, 32'sd793, 32'sd113,
32'sd136, 32'sd324, 32'sd118, 32'sd1189, 32'sd369, 32'sd1978,
32'sd1770, 32'sd345, 32'sd1477, 32'sd257, 32'sd1082, 32'sd647,
32'sd1904, 32'sd1553, 32'sd525, 32'sd512, 32'sd1202, 32'sd995,
32'sd245, 32'sd255, 32'sd1592, 32'sd1324, 32'sd1038, 32'sd664,
32'sd1130, 32'sd1041, 32'sd1487, 32'sd1399, 32'sd138, 32'sd1050,
32'sd1918, 32'sd795, 32'sd1367, 32'sd753, 32'sd269, 32'sd340,
32'sd1381, 32'sd683, 32'sd1549, 32'sd1314, 32'sd1479, 32'sd367,
32'sd477, 32'sd880, 32'sd1392, 32'sd685, 32'sd1841, 32'sd1577,
32'sd1690, 32'sd1670, 32'sd1174, 32'sd1577, 32'sd699, 32'sd497,
32'sd717, 32'sd609, 32'sd1450, 32'sd700, 32'sd1671, 32'sd1167,
32'sd387, 32'sd1962, 32'sd636, 32'sd286, 32'sd1365, 32'sd1459,
32'sd786, 32'sd1696, 32'sd653, 32'sd915, 32'sd1763, 32'sd248,
32'sd1101, 32'sd1993, 32'sd1410, 32'sd1213, 32'sd1701, 32'sd987,
32'sd568, 32'sd620, 32'sd440, 32'sd1354, 32'sd570, 32'sd273,
32'sd795, 32'sd705, 32'sd1808, 32'sd1360, 32'sd1051, 32'sd496,
32'sd1896, 32'sd762, 32'sd1230, 32'sd1726, 32'sd513, 32'sd1495,
32'sd802, 32'sd342, 32'sd1439, 32'sd857, 32'sd303, 32'sd147,
32'sd1130, 32'sd780, 32'sd1325, 32'sd247, 32'sd1842, 32'sd1862,
32'sd469, 32'sd1195, 32'sd1370, 32'sd1463, 32'sd1469, 32'sd725,
32'sd660, 32'sd254, 32'sd469, 32'sd622, 32'sd1077, 32'sd848,
32'sd1197, 32'sd1142, 32'sd1253, 32'sd177, 32'sd1302, 32'sd1547,
32'sd1704, 32'sd742, 32'sd451, 32'sd966, 32'sd1163, 32'sd1067,
32'sd176, 32'sd777, 32'sd955, 32'sd1895, 32'sd807, 32'sd825,
32'sd1448, 32'sd1477, 32'sd1129, 32'sd815, 32'sd1660, 32'sd491,
32'sd1773, 32'sd1858, 32'sd337, 32'sd577, 32'sd723, 32'sd1885,
32'sd1429, 32'sd1177, 32'sd966, 32'sd536, 32'sd681, 32'sd1607,
32'sd1575, 32'sd972, 32'sd1990, 32'sd929, 32'sd260, 32'sd1603,
32'sd1608, 32'sd1154, 32'sd1504, 32'sd329, 32'sd317, 32'sd741,
32'sd485, 32'sd1178, 32'sd1180, 32'sd305, 32'sd1328, 32'sd1878,
32'sd1728, 32'sd505, 32'sd1117, 32'sd1771, 32'sd144, 32'sd1181,
32'sd1528, 32'sd1125, 32'sd681, 32'sd1344, 32'sd1070, 32'sd774,
32'sd1630, 32'sd1486, 32'sd991, 32'sd1174, 32'sd1860, 32'sd1356,
32'sd435, 32'sd748, 32'sd484, 32'sd503, 32'sd437, 32'sd1438,
32'sd161, 32'sd1398, 32'sd773, 32'sd1171, 32'sd591, 32'sd1963,
32'sd1549, 32'sd930, 32'sd116, 32'sd155, 32'sd1223, 32'sd674,
32'sd1244, 32'sd1455, 32'sd223, 32'sd1288, 32'sd1439, 32'sd577,
32'sd1178, 32'sd1897, 32'sd1976, 32'sd1792, 32'sd962, 32'sd1069,
32'sd961, 32'sd1234, 32'sd170, 32'sd1050, 32'sd164, 32'sd1519,
32'sd982, 32'sd1620, 32'sd1712, 32'sd1368, 32'sd1215, 32'sd1609,
32'sd569, 32'sd376, 32'sd1920, 32'sd1518, 32'sd1873, 32'sd1178,
32'sd951, 32'sd1900, 32'sd953, 32'sd1067, 32'sd659, 32'sd862,
32'sd116, 32'sd1387, 32'sd176, 32'sd968, 32'sd1717, 32'sd135,
32'sd1998, 32'sd1970, 32'sd1227, 32'sd432, 32'sd993, 32'sd1172,
32'sd1600, 32'sd1658, 32'sd1022, 32'sd1501, 32'sd773, 32'sd1587,
32'sd194, 32'sd645, 32'sd1985, 32'sd1497, 32'sd1924, 32'sd514,
32'sd398, 32'sd771, 32'sd609, 32'sd1582, 32'sd758, 32'sd1703,
32'sd1162, 32'sd489, 32'sd271, 32'sd1408, 32'sd1483, 32'sd1932,
32'sd122, 32'sd1225, 32'sd981, 32'sd971, 32'sd679, 32'sd396,
32'sd1324, 32'sd1921, 32'sd1980, 32'sd1162, 32'sd375, 32'sd969,
32'sd1286, 32'sd1681, 32'sd924, 32'sd1709, 32'sd1982, 32'sd1215,
32'sd1745, 32'sd913, 32'sd1451, 32'sd638, 32'sd1355, 32'sd1288,
32'sd596, 32'sd1649, 32'sd494, 32'sd1645, 32'sd949, 32'sd566,
32'sd821, 32'sd732, 32'sd665, 32'sd130, 32'sd415, 32'sd465,
32'sd1305, 32'sd918, 32'sd658, 32'sd279, 32'sd1027, 32'sd1399,
32'sd509, 32'sd1167, 32'sd1440, 32'sd676, 32'sd673, 32'sd1080,
32'sd597, 32'sd943, 32'sd1541, 32'sd1297, 32'sd1702, 32'sd323,
32'sd1244, 32'sd559, 32'sd487, 32'sd435, 32'sd533, 32'sd958,
32'sd214, 32'sd174, 32'sd216, 32'sd696, 32'sd984, 32'sd1349,
32'sd1228, 32'sd906, 32'sd174, 32'sd1201, 32'sd543, 32'sd1461,
32'sd387, 32'sd1534, 32'sd1620, 32'sd340, 32'sd267, 32'sd1324,
32'sd223, 32'sd1829, 32'sd292, 32'sd972, 32'sd1077, 32'sd1435,
32'sd169, 32'sd476, 32'sd1894, 32'sd875, 32'sd1987, 32'sd853,
32'sd393, 32'sd386, 32'sd210, 32'sd1850, 32'sd1038, 32'sd456,
32'sd1697, 32'sd1945, 32'sd508, 32'sd150, 32'sd283, 32'sd600,
32'sd711, 32'sd289, 32'sd1650, 32'sd1227, 32'sd784, 32'sd1652,
32'sd758, 32'sd1674, 32'sd1605, 32'sd1323, 32'sd1294, 32'sd1068,
32'sd965, 32'sd1702, 32'sd615, 32'sd938, 32'sd1549, 32'sd241,
32'sd1379, 32'sd568, 32'sd1041, 32'sd941, 32'sd969, 32'sd1526,
32'sd716, 32'sd455, 32'sd1165, 32'sd1710, 32'sd1046, 32'sd1687,
32'sd1065, 32'sd1202, 32'sd1197, 32'sd604, 32'sd1681, 32'sd100,
32'sd1237, 32'sd300, 32'sd1104, 32'sd799, 32'sd1699, 32'sd645,
32'sd397, 32'sd1392, 32'sd1609, 32'sd420, 32'sd1626, 32'sd1007,
32'sd1583, 32'sd1202, 32'sd1358, 32'sd1044, 32'sd157, 32'sd1532,
32'sd809, 32'sd861, 32'sd1185, 32'sd1997, 32'sd896, 32'sd1921,
32'sd1755, 32'sd596, 32'sd1834, 32'sd1452, 32'sd532, 32'sd1460,
32'sd1286, 32'sd1500, 32'sd1190, 32'sd952, 32'sd1218, 32'sd1198,
32'sd1967, 32'sd356, 32'sd288, 32'sd205, 32'sd1883, 32'sd1419,
32'sd495, 32'sd1085, 32'sd1217, 32'sd1186, 32'sd727, 32'sd261,
32'sd458, 32'sd726, 32'sd698, 32'sd515, 32'sd1196, 32'sd1276,
32'sd725, 32'sd1282, 32'sd1259, 32'sd728, 32'sd748, 32'sd466,
32'sd1730, 32'sd1427, 32'sd166, 32'sd668, 32'sd1685, 32'sd1203,
32'sd133, 32'sd909, 32'sd689, 32'sd263, 32'sd109, 32'sd266,
32'sd1512, 32'sd928, 32'sd1021, 32'sd219, 32'sd1083, 32'sd1191,
32'sd337, 32'sd410, 32'sd1558, 32'sd773, 32'sd1233, 32'sd1192,
32'sd1073, 32'sd1279, 32'sd1912, 32'sd671, 32'sd555, 32'sd849,
32'sd668, 32'sd379, 32'sd1910, 32'sd1335, 32'sd1701, 32'sd542,
32'sd1582, 32'sd1471, 32'sd223, 32'sd323, 32'sd1145, 32'sd871,
32'sd240, 32'sd1153, 32'sd1591, 32'sd572, 32'sd1286, 32'sd1425,
32'sd586, 32'sd163, 32'sd1881, 32'sd353, 32'sd790, 32'sd265,
32'sd667, 32'sd333, 32'sd128, 32'sd1115, 32'sd1227, 32'sd802,
32'sd1404, 32'sd327, 32'sd861, 32'sd865, 32'sd138, 32'sd589,
32'sd926, 32'sd575, 32'sd1397, 32'sd1921, 32'sd1052, 32'sd1317,
32'sd892, 32'sd810, 32'sd1737, 32'sd1428, 32'sd1639, 32'sd190,
32'sd917, 32'sd657, 32'sd1941, 32'sd1261, 32'sd166, 32'sd1950,
32'sd1915, 32'sd923, 32'sd221, 32'sd366, 32'sd687, 32'sd591,
32'sd910, 32'sd1164, 32'sd1518, 32'sd729, 32'sd328, 32'sd632,
32'sd706, 32'sd1148, 32'sd1712, 32'sd510, 32'sd129, 32'sd228,
32'sd1857, 32'sd1322, 32'sd844, 32'sd401, 32'sd1375, 32'sd1143,
32'sd1376, 32'sd1848, 32'sd307, 32'sd1694, 32'sd637, 32'sd905,
32'sd731, 32'sd1899, 32'sd1713, 32'sd1252, 32'sd1826, 32'sd215,
32'sd501, 32'sd1985, 32'sd916, 32'sd384, 32'sd1121, 32'sd722,
32'sd158, 32'sd1775, 32'sd693, 32'sd408, 32'sd392, 32'sd1416,
32'sd1009, 32'sd526, 32'sd1842, 32'sd1903, 32'sd236, 32'sd1882,
32'sd1903, 32'sd989, 32'sd1637, 32'sd1781, 32'sd780, 32'sd612,
32'sd1687, 32'sd770, 32'sd558, 32'sd649, 32'sd374, 32'sd370,
32'sd1088, 32'sd1132, 32'sd244, 32'sd777, 32'sd1844, 32'sd1440,
32'sd1884, 32'sd1560, 32'sd453, 32'sd1049, 32'sd529, 32'sd518,
32'sd1524, 32'sd761, 32'sd1406, 32'sd229, 32'sd1014, 32'sd309,
32'sd1960, 32'sd1141, 32'sd1362, 32'sd1236, 32'sd1186, 32'sd1177,
32'sd1232, 32'sd1343, 32'sd546, 32'sd649, 32'sd540, 32'sd1555,
32'sd719, 32'sd863, 32'sd285, 32'sd767, 32'sd1807, 32'sd826,
32'sd649, 32'sd734, 32'sd1407, 32'sd1110, 32'sd1836, 32'sd614,
32'sd192, 32'sd1383, 32'sd307, 32'sd851, 32'sd1616, 32'sd1155,
32'sd1434, 32'sd890, 32'sd612, 32'sd189, 32'sd1743, 32'sd969,
32'sd1156, 32'sd433, 32'sd1540, 32'sd1146, 32'sd130, 32'sd870,
32'sd250, 32'sd384, 32'sd1395, 32'sd1013, 32'sd254, 32'sd392,
32'sd1621, 32'sd1774, 32'sd215, 32'sd242, 32'sd952, 32'sd1884,
32'sd446, 32'sd332, 32'sd125, 32'sd1496, 32'sd815, 32'sd1361,
32'sd1602, 32'sd1227, 32'sd877, 32'sd1114, 32'sd1286, 32'sd107,
32'sd388, 32'sd831, 32'sd1553, 32'sd864, 32'sd243, 32'sd1084,
32'sd1516, 32'sd356, 32'sd1454, 32'sd718, 32'sd1282, 32'sd1216,
32'sd1650, 32'sd273, 32'sd419, 32'sd1752, 32'sd1754, 32'sd1023,
32'sd743, 32'sd624, 32'sd932, 32'sd1110, 32'sd528, 32'sd1457,
32'sd1888, 32'sd1156, 32'sd348, 32'sd1669, 32'sd343, 32'sd477,
32'sd1380, 32'sd540, 32'sd1399, 32'sd681, 32'sd1477, 32'sd1828,
32'sd807, 32'sd1513, 32'sd1004, 32'sd1968, 32'sd147, 32'sd465,
32'sd1884, 32'sd470, 32'sd1272, 32'sd1610, 32'sd1125, 32'sd103,
32'sd259, 32'sd1986, 32'sd316, 32'sd1242, 32'sd1493, 32'sd377,
32'sd515, 32'sd1787, 32'sd899, 32'sd612, 32'sd626, 32'sd479,
32'sd1944, 32'sd1141, 32'sd1686, 32'sd1803, 32'sd1855, 32'sd1579,
32'sd593, 32'sd743, 32'sd1801, 32'sd1625, 32'sd240, 32'sd408,
32'sd1697, 32'sd1803, 32'sd294, 32'sd1968, 32'sd577, 32'sd1030,
32'sd127, 32'sd142, 32'sd1656, 32'sd1269, 32'sd591, 32'sd1524,
32'sd1364, 32'sd376, 32'sd935, 32'sd1329, 32'sd1065, 32'sd563,
32'sd1652, 32'sd430, 32'sd1261, 32'sd1882, 32'sd1372, 32'sd1369,
32'sd1882, 32'sd120, 32'sd908, 32'sd1311, 32'sd1951, 32'sd1704,
32'sd581, 32'sd1004, 32'sd953, 32'sd250, 32'sd832, 32'sd1893,
32'sd261, 32'sd163, 32'sd1099, 32'sd1911, 32'sd1876, 32'sd227,
32'sd838, 32'sd363, 32'sd1156, 32'sd1921, 32'sd856, 32'sd254,
32'sd646, 32'sd1765, 32'sd991, 32'sd1967, 32'sd519, 32'sd549,
32'sd1108, 32'sd216, 32'sd1499, 32'sd859, 32'sd1963, 32'sd669,
32'sd1196, 32'sd1931, 32'sd1878, 32'sd648, 32'sd914, 32'sd1538,
32'sd1503, 32'sd1573, 32'sd1671, 32'sd1052, 32'sd1424, 32'sd1647,
32'sd1206, 32'sd450, 32'sd340, 32'sd458, 32'sd300, 32'sd213,
32'sd1628, 32'sd438, 32'sd389, 32'sd328, 32'sd1631, 32'sd618,
32'sd919, 32'sd507, 32'sd846, 32'sd572, 32'sd618, 32'sd1726,
32'sd1208, 32'sd1627, 32'sd597, 32'sd1550, 32'sd820, 32'sd1392,
32'sd1689, 32'sd1590, 32'sd472, 32'sd1350, 32'sd406, 32'sd1303,
32'sd347, 32'sd862, 32'sd549, 32'sd224, 32'sd1580, 32'sd1513,
32'sd1921, 32'sd1006, 32'sd1525, 32'sd1440, 32'sd1947, 32'sd1536,
32'sd1270, 32'sd1810, 32'sd1240, 32'sd1503, 32'sd969, 32'sd1493,
32'sd1748, 32'sd1057, 32'sd1827, 32'sd1239, 32'sd654, 32'sd222,
32'sd346, 32'sd249, 32'sd1637, 32'sd852, 32'sd691, 32'sd1442,
32'sd1227, 32'sd1880, 32'sd1930, 32'sd1373, 32'sd609, 32'sd149,
32'sd754, 32'sd1362, 32'sd1719, 32'sd750, 32'sd472, 32'sd1835,
32'sd898, 32'sd1452, 32'sd751, 32'sd410, 32'sd442, 32'sd181,
32'sd844, 32'sd1821, 32'sd991, 32'sd1568, 32'sd1101, 32'sd811,
32'sd1636, 32'sd413, 32'sd1718, 32'sd843, 32'sd1551, 32'sd173,
32'sd609, 32'sd785, 32'sd1961, 32'sd553, 32'sd182, 32'sd898,
32'sd1854, 32'sd1968, 32'sd1428, 32'sd1651, 32'sd1576, 32'sd1970,
32'sd766, 32'sd784, 32'sd1252, 32'sd1210, 32'sd1831, 32'sd1324,
32'sd1408, 32'sd466, 32'sd280, 32'sd519, 32'sd1451, 32'sd1640,
32'sd928, 32'sd271, 32'sd513, 32'sd1859, 32'sd1968, 32'sd1586,
32'sd303, 32'sd1898, 32'sd1418, 32'sd1752, 32'sd1950, 32'sd741,
32'sd1082, 32'sd1306, 32'sd1811, 32'sd411, 32'sd1085, 32'sd364,
32'sd806, 32'sd458, 32'sd426, 32'sd1925, 32'sd1945, 32'sd1690,
32'sd1003, 32'sd941, 32'sd317, 32'sd723, 32'sd874, 32'sd1710,
32'sd1668, 32'sd822, 32'sd950, 32'sd205, 32'sd1787, 32'sd1791,
32'sd491, 32'sd828, 32'sd1514, 32'sd579, 32'sd1616, 32'sd1279,
32'sd170, 32'sd1469, 32'sd929, 32'sd1754, 32'sd943, 32'sd495,
32'sd1215, 32'sd1850, 32'sd814, 32'sd1989, 32'sd768, 32'sd799,
32'sd1665, 32'sd1795, 32'sd260, 32'sd625, 32'sd186, 32'sd1241,
32'sd573, 32'sd175, 32'sd347, 32'sd1952, 32'sd1998, 32'sd979,
32'sd947, 32'sd1792, 32'sd808, 32'sd1005, 32'sd697, 32'sd787,
32'sd738, 32'sd688, 32'sd1162, 32'sd1110, 32'sd251, 32'sd1627,
32'sd493, 32'sd1025, 32'sd1279, 32'sd363, 32'sd1771, 32'sd508,
32'sd758, 32'sd952, 32'sd771, 32'sd1744, 32'sd886, 32'sd836,
32'sd1196, 32'sd1527, 32'sd813, 32'sd1816, 32'sd1775, 32'sd1925,
32'sd1718, 32'sd1422, 32'sd1153, 32'sd1514, 32'sd1789, 32'sd1874,
32'sd916, 32'sd1903, 32'sd534, 32'sd746, 32'sd545, 32'sd517,
32'sd813, 32'sd884, 32'sd852, 32'sd1803, 32'sd1369, 32'sd1243,
32'sd833, 32'sd1045, 32'sd479, 32'sd839, 32'sd167, 32'sd355,
32'sd788, 32'sd228, 32'sd766, 32'sd1881, 32'sd1393, 32'sd1209,
32'sd1005, 32'sd921, 32'sd1823, 32'sd970, 32'sd942, 32'sd683,
32'sd411, 32'sd496, 32'sd102, 32'sd1444, 32'sd1732, 32'sd1526,
32'sd471, 32'sd1997, 32'sd513, 32'sd1733, 32'sd1748, 32'sd1588,
32'sd1073, 32'sd619, 32'sd1048, 32'sd1251, 32'sd1264, 32'sd1734,
32'sd205, 32'sd1697, 32'sd1026, 32'sd1700, 32'sd293, 32'sd930,
32'sd707, 32'sd1834, 32'sd1427, 32'sd1005, 32'sd674, 32'sd1161,
32'sd980, 32'sd1453, 32'sd313, 32'sd1304, 32'sd134, 32'sd1985,
32'sd1913, 32'sd462, 32'sd884, 32'sd794, 32'sd1537, 32'sd1940,
32'sd1248, 32'sd1657, 32'sd228, 32'sd1917, 32'sd978, 32'sd409,
32'sd350, 32'sd1477, 32'sd1282, 32'sd1181, 32'sd1136, 32'sd1478,
32'sd1117, 32'sd1391, 32'sd604, 32'sd1017, 32'sd348, 32'sd273,
32'sd1748, 32'sd443, 32'sd1702, 32'sd642, 32'sd568, 32'sd1227,
32'sd1872, 32'sd679, 32'sd1108, 32'sd1050, 32'sd1120, 32'sd387,
32'sd1055, 32'sd1456, 32'sd481, 32'sd1761, 32'sd1975, 32'sd774,
32'sd1707, 32'sd701, 32'sd882, 32'sd1762, 32'sd610, 32'sd757,
32'sd1869, 32'sd1172, 32'sd1109, 32'sd784, 32'sd1687, 32'sd1790,
32'sd1185, 32'sd931, 32'sd1196, 32'sd722, 32'sd1418, 32'sd647,
32'sd1363, 32'sd308, 32'sd1051, 32'sd130, 32'sd911, 32'sd1062,
32'sd132, 32'sd1397, 32'sd636, 32'sd296, 32'sd934, 32'sd620,
32'sd294, 32'sd1725, 32'sd1311, 32'sd1257, 32'sd632, 32'sd1474,
32'sd1324, 32'sd1002, 32'sd1636, 32'sd1029, 32'sd1058, 32'sd1837,
32'sd315, 32'sd904, 32'sd1125, 32'sd1595, 32'sd1791, 32'sd1281,
32'sd505, 32'sd455, 32'sd665, 32'sd1950, 32'sd916, 32'sd1269,
32'sd435, 32'sd759, 32'sd263, 32'sd458, 32'sd109, 32'sd1736,
32'sd1864, 32'sd1945, 32'sd862, 32'sd1933, 32'sd502, 32'sd1250,
32'sd713, 32'sd1133, 32'sd1104, 32'sd907, 32'sd394, 32'sd419,
32'sd598, 32'sd204, 32'sd968, 32'sd899, 32'sd1527, 32'sd779,
32'sd1678, 32'sd710, 32'sd1364, 32'sd1339, 32'sd1737, 32'sd652,
32'sd171, 32'sd645, 32'sd1831, 32'sd988, 32'sd1780, 32'sd1576,
32'sd903, 32'sd1431, 32'sd1082, 32'sd464, 32'sd1836, 32'sd1144,
32'sd1086, 32'sd1201, 32'sd679, 32'sd1341, 32'sd648, 32'sd532,
32'sd1294, 32'sd1860, 32'sd1056, 32'sd1794, 32'sd811, 32'sd982,
32'sd950, 32'sd846, 32'sd244, 32'sd608, 32'sd795, 32'sd110,
32'sd982, 32'sd716, 32'sd1040, 32'sd1756, 32'sd589, 32'sd1512,
32'sd345, 32'sd1164, 32'sd741, 32'sd425, 32'sd908, 32'sd290,
32'sd1592, 32'sd1189, 32'sd1068, 32'sd565, 32'sd1059, 32'sd1495,
32'sd1414, 32'sd1238, 32'sd1181, 32'sd334, 32'sd1606, 32'sd1378,
32'sd1217, 32'sd1866, 32'sd1215, 32'sd807, 32'sd1106, 32'sd701,
32'sd1416, 32'sd896, 32'sd1713, 32'sd109, 32'sd1017, 32'sd1674,
32'sd1453, 32'sd1220, 32'sd364, 32'sd233, 32'sd1904, 32'sd416,
32'sd777, 32'sd767, 32'sd1479, 32'sd347, 32'sd1939, 32'sd1402,
32'sd204, 32'sd343, 32'sd928, 32'sd187, 32'sd680, 32'sd682,
32'sd1493, 32'sd608, 32'sd734, 32'sd1746, 32'sd266, 32'sd618,
32'sd1403, 32'sd1006, 32'sd260, 32'sd474, 32'sd1965, 32'sd463,
32'sd1852, 32'sd1016, 32'sd1780, 32'sd210, 32'sd1982, 32'sd306,
32'sd1827, 32'sd277, 32'sd118, 32'sd1061, 32'sd451, 32'sd1183,
32'sd1397, 32'sd1257, 32'sd438, 32'sd1289, 32'sd583, 32'sd1895,
32'sd510, 32'sd269, 32'sd1280, 32'sd421, 32'sd1391, 32'sd1209,
32'sd847, 32'sd1679, 32'sd1770, 32'sd1969, 32'sd383, 32'sd301,
32'sd1841, 32'sd134, 32'sd1109, 32'sd653, 32'sd952, 32'sd1877,
32'sd106, 32'sd1444, 32'sd1876, 32'sd1347, 32'sd1846, 32'sd203,
32'sd1878, 32'sd375, 32'sd663, 32'sd1620, 32'sd1079, 32'sd606,
32'sd1943, 32'sd968, 32'sd1820, 32'sd357, 32'sd1607, 32'sd296,
32'sd601, 32'sd1131, 32'sd168, 32'sd867, 32'sd1265, 32'sd528,
32'sd779, 32'sd401, 32'sd1053, 32'sd1412, 32'sd1401, 32'sd1188,
32'sd1364, 32'sd239, 32'sd983, 32'sd667, 32'sd946, 32'sd1431,
32'sd1428, 32'sd1621, 32'sd434, 32'sd945, 32'sd918, 32'sd1497,
32'sd892, 32'sd383, 32'sd782, 32'sd793, 32'sd1166, 32'sd697,
32'sd841, 32'sd1584, 32'sd200, 32'sd1062, 32'sd223, 32'sd732,
32'sd1895, 32'sd1168, 32'sd559, 32'sd1640, 32'sd920, 32'sd803,
32'sd679, 32'sd1141, 32'sd1253, 32'sd1286, 32'sd321, 32'sd488,
32'sd569, 32'sd1437, 32'sd1212, 32'sd1652, 32'sd221, 32'sd930,
32'sd948, 32'sd1217, 32'sd1662, 32'sd119, 32'sd170, 32'sd839,
32'sd889, 32'sd727, 32'sd445, 32'sd1733, 32'sd1611, 32'sd164,
32'sd306, 32'sd786, 32'sd1490, 32'sd1316, 32'sd105, 32'sd192,
32'sd1328, 32'sd1735, 32'sd1005, 32'sd575, 32'sd742, 32'sd1028,
32'sd362, 32'sd1156, 32'sd516, 32'sd764, 32'sd1821, 32'sd1001,
32'sd1002, 32'sd1717, 32'sd456, 32'sd537, 32'sd1361, 32'sd116,
32'sd127, 32'sd1251, 32'sd1375, 32'sd969, 32'sd1138, 32'sd1346,
32'sd1119, 32'sd697, 32'sd392, 32'sd1028, 32'sd1916, 32'sd785,
32'sd195, 32'sd481, 32'sd152, 32'sd1004, 32'sd1163, 32'sd1058,
32'sd787, 32'sd438, 32'sd1834, 32'sd1061, 32'sd1956, 32'sd513,
32'sd641, 32'sd1096, 32'sd1493, 32'sd1614, 32'sd1204, 32'sd1613,
32'sd1158, 32'sd1302, 32'sd1397, 32'sd1045, 32'sd275, 32'sd492,
32'sd578, 32'sd811, 32'sd1273, 32'sd1930, 32'sd1361, 32'sd1730,
32'sd732, 32'sd201, 32'sd785, 32'sd1524, 32'sd1357, 32'sd1420,
32'sd571, 32'sd1756, 32'sd174, 32'sd840, 32'sd857, 32'sd1764,
32'sd1444, 32'sd469, 32'sd928, 32'sd299, 32'sd1203, 32'sd1960,
32'sd1271, 32'sd1401, 32'sd1932, 32'sd331, 32'sd1280, 32'sd1318,
32'sd985, 32'sd598, 32'sd632, 32'sd1962, 32'sd830, 32'sd1928,
32'sd636, 32'sd225, 32'sd261, 32'sd613, 32'sd1983, 32'sd535,
32'sd721, 32'sd1257, 32'sd1325, 32'sd1958, 32'sd1351, 32'sd1663,
32'sd1657, 32'sd1941, 32'sd545, 32'sd1606, 32'sd916, 32'sd191,
32'sd1177, 32'sd1097, 32'sd1254, 32'sd235, 32'sd1025, 32'sd823,
32'sd1842, 32'sd1663, 32'sd314, 32'sd914, 32'sd1718, 32'sd1920,
32'sd731, 32'sd797, 32'sd330, 32'sd1106, 32'sd317, 32'sd300,
32'sd1216, 32'sd1675, 32'sd780, 32'sd161, 32'sd570, 32'sd1503,
32'sd1970, 32'sd779, 32'sd1391, 32'sd1477, 32'sd1609, 32'sd1313,
32'sd371, 32'sd754, 32'sd1357, 32'sd205, 32'sd843, 32'sd1319,
32'sd1370, 32'sd185, 32'sd1740, 32'sd1815, 32'sd412, 32'sd522,
32'sd1865, 32'sd764, 32'sd1288, 32'sd1120, 32'sd620, 32'sd1419,
32'sd766, 32'sd1804, 32'sd813, 32'sd184, 32'sd1228, 32'sd1287,
32'sd1016, 32'sd1455, 32'sd204, 32'sd1672, 32'sd446, 32'sd689,
32'sd1604, 32'sd1105, 32'sd1740, 32'sd337, 32'sd1205, 32'sd475,
32'sd1492, 32'sd222, 32'sd967, 32'sd1320, 32'sd310, 32'sd1307,
32'sd837, 32'sd1013, 32'sd1997, 32'sd267, 32'sd1216, 32'sd300,
32'sd561, 32'sd1901, 32'sd552, 32'sd1214, 32'sd1751, 32'sd1533,
32'sd1261, 32'sd1742, 32'sd1249, 32'sd415, 32'sd149, 32'sd1727,
32'sd1296, 32'sd883, 32'sd958, 32'sd1590, 32'sd165, 32'sd1951,
32'sd124, 32'sd1155, 32'sd1576, 32'sd161, 32'sd687, 32'sd443,
32'sd1905, 32'sd561, 32'sd1424, 32'sd441, 32'sd1082, 32'sd762,
32'sd1038, 32'sd1118, 32'sd1001, 32'sd487, 32'sd1966, 32'sd218,
32'sd1198, 32'sd170, 32'sd639, 32'sd318, 32'sd226, 32'sd1441,
32'sd1365, 32'sd807, 32'sd557, 32'sd406, 32'sd284, 32'sd1242,
32'sd112, 32'sd1896, 32'sd148, 32'sd432, 32'sd112, 32'sd671,
32'sd1675, 32'sd701, 32'sd1939, 32'sd301, 32'sd884, 32'sd167,
32'sd428, 32'sd296, 32'sd1532, 32'sd901, 32'sd1345, 32'sd544,
32'sd1290, 32'sd932, 32'sd1078, 32'sd1290, 32'sd1064, 32'sd733,
32'sd591, 32'sd915, 32'sd1281, 32'sd721, 32'sd1380, 32'sd1537,
32'sd635, 32'sd1159, 32'sd1972, 32'sd571, 32'sd1850, 32'sd1080,
32'sd1062, 32'sd421, 32'sd1492, 32'sd1397, 32'sd1635, 32'sd180,
32'sd438, 32'sd448, 32'sd1204, 32'sd1771, 32'sd399, 32'sd1039,
32'sd922, 32'sd762, 32'sd1033, 32'sd629, 32'sd1710, 32'sd1024,
32'sd1329, 32'sd1366, 32'sd1176, 32'sd1405, 32'sd1049, 32'sd530,
32'sd1412, 32'sd1868, 32'sd353, 32'sd1795, 32'sd272, 32'sd1347,
32'sd592, 32'sd956, 32'sd1717, 32'sd1364, 32'sd1390, 32'sd233,
32'sd578, 32'sd913, 32'sd1655, 32'sd1726, 32'sd1419, 32'sd1590,
32'sd846, 32'sd935, 32'sd435, 32'sd193, 32'sd696, 32'sd1040,
32'sd1212, 32'sd1884, 32'sd909, 32'sd670, 32'sd1318, 32'sd571,
32'sd463, 32'sd853, 32'sd1834, 32'sd326, 32'sd1787, 32'sd549,
32'sd1223, 32'sd1318, 32'sd523, 32'sd1180, 32'sd1416, 32'sd994,
32'sd1316, 32'sd343, 32'sd1901, 32'sd1855, 32'sd1133, 32'sd1586,
32'sd1994, 32'sd202, 32'sd936, 32'sd1823, 32'sd1153, 32'sd1038,
32'sd399, 32'sd751, 32'sd1292, 32'sd629, 32'sd135, 32'sd408,
32'sd1890, 32'sd1050, 32'sd1551, 32'sd1855, 32'sd1966, 32'sd884,
32'sd258, 32'sd1411, 32'sd324, 32'sd1593, 32'sd1512, 32'sd1073,
32'sd392, 32'sd1350, 32'sd1785, 32'sd1673, 32'sd663, 32'sd1356,
32'sd1169, 32'sd127, 32'sd115, 32'sd1000, 32'sd1558, 32'sd243,
32'sd1213, 32'sd1221, 32'sd855, 32'sd534, 32'sd588, 32'sd1558,
32'sd968, 32'sd396, 32'sd627, 32'sd956, 32'sd849, 32'sd1293,
32'sd503, 32'sd751, 32'sd661, 32'sd1545, 32'sd1339, 32'sd1742,
32'sd1006, 32'sd725, 32'sd480, 32'sd160, 32'sd1658, 32'sd172,
32'sd1344, 32'sd408, 32'sd164, 32'sd307, 32'sd1809, 32'sd1857,
32'sd1392, 32'sd300, 32'sd973, 32'sd856, 32'sd181, 32'sd940,
32'sd679, 32'sd936, 32'sd1666, 32'sd1090, 32'sd830, 32'sd1701,
32'sd1788, 32'sd426, 32'sd1488, 32'sd1100, 32'sd709, 32'sd774,
32'sd1749, 32'sd1340, 32'sd524, 32'sd885, 32'sd1023, 32'sd265,
32'sd1366, 32'sd1622, 32'sd374, 32'sd280, 32'sd327, 32'sd1415,
32'sd1292, 32'sd1403, 32'sd1570, 32'sd111, 32'sd1571, 32'sd1058,
32'sd1075, 32'sd1209, 32'sd782, 32'sd1664, 32'sd1222, 32'sd369,
32'sd320, 32'sd1064, 32'sd413, 32'sd1946, 32'sd991, 32'sd1704,
32'sd1470, 32'sd558, 32'sd1007, 32'sd754, 32'sd1079, 32'sd975,
32'sd659, 32'sd1724, 32'sd1994, 32'sd1205, 32'sd529, 32'sd807,
32'sd1170, 32'sd376, 32'sd1640, 32'sd1274, 32'sd797, 32'sd1691,
32'sd858, 32'sd1124, 32'sd1531, 32'sd535, 32'sd598, 32'sd423,
32'sd1052, 32'sd1891, 32'sd622, 32'sd1369, 32'sd955, 32'sd1929,
32'sd311, 32'sd341, 32'sd294, 32'sd544, 32'sd358, 32'sd1802,
32'sd861, 32'sd1340, 32'sd1416, 32'sd1895, 32'sd1085, 32'sd1813,
32'sd978, 32'sd1890, 32'sd1968, 32'sd888, 32'sd1358, 32'sd683,
32'sd793, 32'sd1069, 32'sd1453, 32'sd192, 32'sd320, 32'sd1024,
32'sd1221, 32'sd1067, 32'sd100, 32'sd882, 32'sd1824, 32'sd943,
32'sd1094, 32'sd934, 32'sd704, 32'sd1352, 32'sd626, 32'sd1142,
32'sd823, 32'sd1491, 32'sd1972, 32'sd900, 32'sd331, 32'sd554,
32'sd1725, 32'sd1189, 32'sd1876, 32'sd742, 32'sd1388, 32'sd856,
32'sd116, 32'sd1164, 32'sd734, 32'sd1591, 32'sd1154, 32'sd1399,
32'sd1143, 32'sd542, 32'sd1541, 32'sd334, 32'sd943, 32'sd1964,
32'sd1853, 32'sd1012, 32'sd1590, 32'sd771, 32'sd1239, 32'sd1363,
32'sd1151, 32'sd1972, 32'sd474, 32'sd1957, 32'sd344, 32'sd1915,
32'sd599, 32'sd306, 32'sd1969, 32'sd1999, 32'sd802, 32'sd213,
32'sd1173, 32'sd1104, 32'sd739, 32'sd480, 32'sd636, 32'sd903,
32'sd754, 32'sd882, 32'sd104, 32'sd1011, 32'sd921, 32'sd831,
32'sd260, 32'sd321, 32'sd550, 32'sd360, 32'sd1403, 32'sd1538,
32'sd396, 32'sd1514, 32'sd1979, 32'sd1257, 32'sd1249, 32'sd843,
32'sd1609, 32'sd211, 32'sd504, 32'sd132, 32'sd1440, 32'sd953,
32'sd1776, 32'sd606, 32'sd1135, 32'sd473, 32'sd1891, 32'sd606,
32'sd811, 32'sd482, 32'sd1965, 32'sd1100, 32'sd1814, 32'sd1399,
32'sd299, 32'sd1579, 32'sd1783, 32'sd1569, 32'sd1168, 32'sd1026,
32'sd345, 32'sd945, 32'sd1656, 32'sd319, 32'sd343, 32'sd350,
32'sd348, 32'sd228, 32'sd341, 32'sd340, 32'sd530, 32'sd781,
32'sd1131, 32'sd1533, 32'sd743, 32'sd873, 32'sd755, 32'sd850,
32'sd621, 32'sd636, 32'sd503, 32'sd1430, 32'sd1589, 32'sd394,
32'sd950, 32'sd1693, 32'sd1876, 32'sd1701, 32'sd318, 32'sd261,
32'sd1264, 32'sd584, 32'sd1060, 32'sd1029, 32'sd1561, 32'sd1548,
32'sd1681, 32'sd737, 32'sd1877, 32'sd228, 32'sd526, 32'sd1881,
32'sd1877, 32'sd143, 32'sd1949, 32'sd769, 32'sd1425, 32'sd952,
32'sd1834, 32'sd426, 32'sd817, 32'sd1794, 32'sd1479, 32'sd1503,
32'sd1308, 32'sd1623, 32'sd267, 32'sd1422, 32'sd788, 32'sd1810,
32'sd609, 32'sd1710, 32'sd1413, 32'sd1948, 32'sd1149, 32'sd576,
32'sd745, 32'sd778, 32'sd1224, 32'sd876, 32'sd1616, 32'sd409,
32'sd623, 32'sd684, 32'sd453, 32'sd1150, 32'sd1379, 32'sd253,
32'sd116, 32'sd1839, 32'sd1951, 32'sd981, 32'sd350, 32'sd1018,
32'sd1254, 32'sd870, 32'sd561, 32'sd779, 32'sd961, 32'sd133,
32'sd1118, 32'sd1752, 32'sd1119, 32'sd199, 32'sd130, 32'sd323,
32'sd929, 32'sd172, 32'sd138, 32'sd1432, 32'sd1769, 32'sd157,
32'sd1429, 32'sd1742, 32'sd1934, 32'sd710, 32'sd1451, 32'sd159,
32'sd937, 32'sd1384, 32'sd289, 32'sd198, 32'sd456, 32'sd1774,
32'sd1626, 32'sd370, 32'sd1241, 32'sd1142, 32'sd336, 32'sd1395,
32'sd1892, 32'sd208, 32'sd533, 32'sd742, 32'sd468, 32'sd1901,
32'sd1928, 32'sd237, 32'sd197, 32'sd1055, 32'sd428, 32'sd228,
32'sd888, 32'sd1979, 32'sd421, 32'sd158, 32'sd833, 32'sd952,
32'sd1345, 32'sd724, 32'sd1715, 32'sd110, 32'sd618, 32'sd1149,
32'sd747, 32'sd344, 32'sd648, 32'sd1368, 32'sd823, 32'sd1183,
32'sd1881, 32'sd600, 32'sd1659, 32'sd810, 32'sd423, 32'sd623,
32'sd1595, 32'sd904, 32'sd784, 32'sd1205, 32'sd986, 32'sd1815,
32'sd1904, 32'sd653, 32'sd191, 32'sd1343, 32'sd535, 32'sd1998,
32'sd1526, 32'sd1815, 32'sd1219, 32'sd568, 32'sd481, 32'sd1785,
32'sd181, 32'sd1541, 32'sd872, 32'sd1038, 32'sd242, 32'sd944,
32'sd1937, 32'sd388, 32'sd759, 32'sd437, 32'sd453, 32'sd483,
32'sd387, 32'sd1941, 32'sd498, 32'sd169, 32'sd376, 32'sd900,
32'sd760, 32'sd1865, 32'sd154, 32'sd123, 32'sd466, 32'sd125,
32'sd193, 32'sd1517, 32'sd1512, 32'sd610, 32'sd1550, 32'sd244,
32'sd1519, 32'sd151, 32'sd1534, 32'sd1703, 32'sd1865, 32'sd816,
32'sd1569, 32'sd1475, 32'sd811, 32'sd1306, 32'sd192, 32'sd1803,
32'sd1338, 32'sd1156, 32'sd882, 32'sd1171, 32'sd589, 32'sd731,
32'sd1820, 32'sd742, 32'sd624, 32'sd180, 32'sd591, 32'sd1184,
32'sd903, 32'sd757, 32'sd1269, 32'sd724, 32'sd559, 32'sd1930,
32'sd1567, 32'sd314, 32'sd702, 32'sd1708, 32'sd1658, 32'sd1474,
32'sd565, 32'sd1211, 32'sd1716, 32'sd948, 32'sd354, 32'sd456,
32'sd1713, 32'sd260, 32'sd1771, 32'sd738, 32'sd968, 32'sd1639,
32'sd1733, 32'sd1860, 32'sd141, 32'sd1334, 32'sd1361, 32'sd1759,
32'sd900, 32'sd290, 32'sd105, 32'sd389, 32'sd793, 32'sd1768,
32'sd1478, 32'sd1295, 32'sd567, 32'sd1584, 32'sd1723, 32'sd1592,
32'sd168, 32'sd250, 32'sd1868, 32'sd1751, 32'sd1313, 32'sd1266,
32'sd917, 32'sd709, 32'sd1474, 32'sd1121, 32'sd1712, 32'sd602,
32'sd1437, 32'sd1504, 32'sd1415, 32'sd1124, 32'sd462, 32'sd726,
32'sd540, 32'sd1520, 32'sd1551, 32'sd1562, 32'sd1462, 32'sd844,
32'sd1291, 32'sd126, 32'sd960, 32'sd213, 32'sd703, 32'sd428,
32'sd1281, 32'sd1002, 32'sd1143, 32'sd1596, 32'sd331, 32'sd1673,
32'sd1438, 32'sd1173, 32'sd871, 32'sd1745, 32'sd345, 32'sd180,
32'sd1337, 32'sd1419, 32'sd907, 32'sd1031, 32'sd620, 32'sd899,
32'sd1777, 32'sd1446, 32'sd992, 32'sd1687, 32'sd1683, 32'sd1194,
32'sd1117, 32'sd727, 32'sd551, 32'sd334, 32'sd218, 32'sd197,
32'sd803, 32'sd1037, 32'sd1358, 32'sd219, 32'sd1063, 32'sd1765,
32'sd1096, 32'sd224, 32'sd180, 32'sd934, 32'sd1933, 32'sd847,
32'sd1541, 32'sd1669, 32'sd1870, 32'sd1187, 32'sd175, 32'sd260,
32'sd1165, 32'sd351, 32'sd1604, 32'sd1061, 32'sd493, 32'sd901,
32'sd1021, 32'sd1862, 32'sd668, 32'sd1876, 32'sd169, 32'sd132,
32'sd1675, 32'sd1867, 32'sd1211, 32'sd1525, 32'sd964, 32'sd450,
32'sd1361, 32'sd1017, 32'sd1876, 32'sd1424, 32'sd500, 32'sd465,
32'sd287, 32'sd530, 32'sd124, 32'sd931, 32'sd212, 32'sd1159,
32'sd1839, 32'sd1312, 32'sd1006, 32'sd702, 32'sd559, 32'sd683,
32'sd1781, 32'sd959, 32'sd1396, 32'sd1126, 32'sd1266, 32'sd383,
32'sd1186, 32'sd1170, 32'sd1857, 32'sd100, 32'sd1649, 32'sd764,
32'sd112, 32'sd1165, 32'sd626, 32'sd871, 32'sd1267, 32'sd174,
32'sd1348, 32'sd738, 32'sd297, 32'sd1852, 32'sd1845, 32'sd1106,
32'sd466, 32'sd1476, 32'sd1996, 32'sd974, 32'sd737, 32'sd286,
32'sd1443, 32'sd243, 32'sd1691, 32'sd777, 32'sd704, 32'sd1013,
32'sd1454, 32'sd1039, 32'sd1582, 32'sd1022, 32'sd1797, 32'sd1821,
32'sd1362, 32'sd1493, 32'sd557, 32'sd1464, 32'sd1250, 32'sd1835,
32'sd667, 32'sd1669, 32'sd1991, 32'sd128, 32'sd1112, 32'sd785,
32'sd106, 32'sd1628, 32'sd205, 32'sd1972, 32'sd866, 32'sd1662,
32'sd558, 32'sd257, 32'sd436, 32'sd344, 32'sd559, 32'sd733,
32'sd1231, 32'sd1357, 32'sd1345, 32'sd1078, 32'sd568, 32'sd1126,
32'sd283, 32'sd1448, 32'sd1204, 32'sd1303, 32'sd896, 32'sd1026,
32'sd1407, 32'sd439, 32'sd940, 32'sd1979, 32'sd391, 32'sd1578,
32'sd1399, 32'sd1776, 32'sd222, 32'sd1329, 32'sd1294, 32'sd477,
32'sd1082, 32'sd1647, 32'sd802, 32'sd146, 32'sd1407, 32'sd1910,
32'sd1084, 32'sd595, 32'sd680, 32'sd898, 32'sd1748, 32'sd895,
32'sd922, 32'sd452, 32'sd832, 32'sd1934, 32'sd664, 32'sd1217,
32'sd1066, 32'sd238, 32'sd1645, 32'sd1300, 32'sd1017, 32'sd1239,
32'sd988, 32'sd633, 32'sd1595, 32'sd1378, 32'sd209, 32'sd1895,
32'sd1924, 32'sd1364, 32'sd809, 32'sd707, 32'sd1571, 32'sd902,
32'sd1692, 32'sd118, 32'sd197, 32'sd678, 32'sd1060, 32'sd1361,
32'sd1418, 32'sd188, 32'sd1385, 32'sd1777, 32'sd415, 32'sd248,
32'sd167, 32'sd1676, 32'sd882, 32'sd891, 32'sd153, 32'sd1139,
32'sd1118, 32'sd1203, 32'sd461, 32'sd544, 32'sd1762, 32'sd1451,
32'sd524, 32'sd1239, 32'sd574, 32'sd1076, 32'sd1086, 32'sd1991,
32'sd422, 32'sd462, 32'sd465, 32'sd1720, 32'sd1990, 32'sd234,
32'sd1530, 32'sd707, 32'sd901, 32'sd1663, 32'sd1090, 32'sd1638,
32'sd1330, 32'sd719, 32'sd1921, 32'sd1101, 32'sd1717, 32'sd1692,
32'sd226, 32'sd769, 32'sd1990, 32'sd562, 32'sd1699, 32'sd1330,
32'sd1977, 32'sd1377, 32'sd457, 32'sd704, 32'sd1917, 32'sd427,
32'sd1800, 32'sd266, 32'sd813, 32'sd1197, 32'sd781, 32'sd1973,
32'sd614, 32'sd715, 32'sd838, 32'sd1234, 32'sd1320, 32'sd552,
32'sd440, 32'sd857, 32'sd1722, 32'sd1888, 32'sd890, 32'sd1543,
32'sd1392, 32'sd1959, 32'sd1065, 32'sd539, 32'sd1557, 32'sd1819,
32'sd1303, 32'sd787, 32'sd1461, 32'sd1923, 32'sd1035, 32'sd1350,
32'sd1312, 32'sd715, 32'sd109, 32'sd924, 32'sd494, 32'sd202,
32'sd1179, 32'sd870, 32'sd1578, 32'sd1859, 32'sd1306, 32'sd1750,
32'sd287, 32'sd1447, 32'sd1945, 32'sd184, 32'sd689, 32'sd957,
32'sd1515, 32'sd1834, 32'sd114, 32'sd462, 32'sd742, 32'sd364,
32'sd192, 32'sd1843, 32'sd1501, 32'sd680, 32'sd1045, 32'sd1331,
32'sd1137, 32'sd1125, 32'sd165, 32'sd281, 32'sd1277, 32'sd1062,
32'sd188, 32'sd1157, 32'sd137, 32'sd778, 32'sd971, 32'sd265,
32'sd152, 32'sd357, 32'sd1540, 32'sd943, 32'sd1399, 32'sd814,
32'sd154, 32'sd1778, 32'sd666, 32'sd1167, 32'sd1032, 32'sd1883,
32'sd1271, 32'sd1163, 32'sd984, 32'sd832, 32'sd780, 32'sd1809,
32'sd1566, 32'sd1820, 32'sd1397, 32'sd275, 32'sd209, 32'sd1584,
32'sd1318, 32'sd591, 32'sd1621, 32'sd1938, 32'sd744, 32'sd896,
32'sd1274, 32'sd1114, 32'sd1304, 32'sd1255, 32'sd1344, 32'sd849,
32'sd1747, 32'sd944, 32'sd1157, 32'sd305, 32'sd1176, 32'sd1686,
32'sd204, 32'sd777, 32'sd1602, 32'sd433, 32'sd241, 32'sd943,
32'sd1260, 32'sd1737, 32'sd281, 32'sd462, 32'sd238, 32'sd1591,
32'sd1949, 32'sd840, 32'sd1960, 32'sd332, 32'sd1633, 32'sd1731,
32'sd511, 32'sd1430, 32'sd814, 32'sd1691, 32'sd1494, 32'sd427,
32'sd398, 32'sd1893, 32'sd403, 32'sd1472, 32'sd373, 32'sd1254,
32'sd1332, 32'sd789, 32'sd292, 32'sd1402, 32'sd1522, 32'sd776,
32'sd524, 32'sd1956, 32'sd103, 32'sd272, 32'sd1323, 32'sd1223,
32'sd1619, 32'sd1765, 32'sd303, 32'sd339, 32'sd1759, 32'sd1359,
32'sd313, 32'sd1023, 32'sd1858, 32'sd1030, 32'sd1279, 32'sd1755,
32'sd261, 32'sd1909, 32'sd1403, 32'sd1585, 32'sd1494, 32'sd803,
32'sd1254, 32'sd1674, 32'sd1980, 32'sd385, 32'sd1499, 32'sd992,
32'sd983, 32'sd956, 32'sd1360, 32'sd1780, 32'sd442, 32'sd1457,
32'sd327, 32'sd1523, 32'sd273, 32'sd1225, 32'sd268, 32'sd1277,
32'sd1087, 32'sd1480, 32'sd764, 32'sd267, 32'sd1173, 32'sd339,
32'sd1731, 32'sd1675, 32'sd1254, 32'sd1494, 32'sd468, 32'sd603,
32'sd1080, 32'sd828, 32'sd515, 32'sd1653, 32'sd953, 32'sd1129,
32'sd884, 32'sd1306, 32'sd633, 32'sd888, 32'sd1198, 32'sd786,
32'sd1325, 32'sd166, 32'sd1397, 32'sd1647, 32'sd762, 32'sd431,
32'sd176, 32'sd1339, 32'sd364, 32'sd667, 32'sd323, 32'sd1855,
32'sd574, 32'sd1837, 32'sd245, 32'sd1895, 32'sd193, 32'sd1345,
32'sd1374, 32'sd1646, 32'sd1575, 32'sd1582, 32'sd1545, 32'sd265,
32'sd1407, 32'sd1963, 32'sd1990, 32'sd1412, 32'sd1432, 32'sd1930,
32'sd1050, 32'sd1775, 32'sd1319, 32'sd1020, 32'sd1752, 32'sd798,
32'sd1959, 32'sd340, 32'sd300, 32'sd237, 32'sd1224, 32'sd1784,
32'sd1585, 32'sd472, 32'sd244, 32'sd869, 32'sd1818, 32'sd967,
32'sd429, 32'sd248, 32'sd513, 32'sd1212, 32'sd115, 32'sd935,
32'sd411, 32'sd1715, 32'sd460, 32'sd1756, 32'sd1773, 32'sd570,
32'sd1770, 32'sd1045, 32'sd1520, 32'sd255, 32'sd658, 32'sd636,
32'sd1160, 32'sd532, 32'sd1612, 32'sd1592, 32'sd1570, 32'sd1750,
32'sd1348, 32'sd1892, 32'sd1141, 32'sd438, 32'sd1697, 32'sd1556,
32'sd1419, 32'sd577, 32'sd729, 32'sd1307, 32'sd110, 32'sd1634,
32'sd1936, 32'sd818, 32'sd1352, 32'sd583, 32'sd1245, 32'sd826,
32'sd305, 32'sd680, 32'sd415, 32'sd489, 32'sd1806, 32'sd890,
32'sd1733, 32'sd652, 32'sd343, 32'sd384, 32'sd743, 32'sd520,
32'sd527, 32'sd579, 32'sd893, 32'sd852, 32'sd1899, 32'sd764,
32'sd524, 32'sd1398, 32'sd948, 32'sd849, 32'sd1315, 32'sd499,
32'sd706, 32'sd1995, 32'sd565, 32'sd1419, 32'sd1167, 32'sd1569,
32'sd144, 32'sd1229, 32'sd121, 32'sd1511, 32'sd1166, 32'sd1632,
32'sd1115, 32'sd703, 32'sd1547, 32'sd1409, 32'sd1446, 32'sd1403,
32'sd1600, 32'sd201, 32'sd916, 32'sd432, 32'sd641, 32'sd1419,
32'sd1325, 32'sd1779, 32'sd1738, 32'sd437, 32'sd509, 32'sd1620,
32'sd878, 32'sd1744, 32'sd1579, 32'sd1168, 32'sd1704, 32'sd1468,
32'sd1553, 32'sd1227, 32'sd615, 32'sd1982, 32'sd1482, 32'sd1109,
32'sd1602, 32'sd1023, 32'sd1344, 32'sd1026, 32'sd1160, 32'sd358,
32'sd554, 32'sd1873, 32'sd1168, 32'sd945, 32'sd674, 32'sd1255,
32'sd366, 32'sd1185, 32'sd1127, 32'sd759, 32'sd616, 32'sd983,
32'sd1371, 32'sd1515, 32'sd1500, 32'sd1684, 32'sd372, 32'sd385,
32'sd107, 32'sd1083, 32'sd1544, 32'sd1771, 32'sd1072, 32'sd216,
32'sd1550, 32'sd1983, 32'sd1962, 32'sd1791, 32'sd1841, 32'sd1073,
32'sd709, 32'sd220, 32'sd1886, 32'sd174, 32'sd179, 32'sd893,
32'sd1361, 32'sd1866, 32'sd383, 32'sd1060, 32'sd1141, 32'sd1534,
32'sd1719, 32'sd1150, 32'sd1935, 32'sd148, 32'sd1537, 32'sd665,
32'sd1089, 32'sd795, 32'sd211, 32'sd1360, 32'sd285, 32'sd1459,
32'sd440, 32'sd1063, 32'sd1801, 32'sd1765, 32'sd1951, 32'sd451,
32'sd709, 32'sd1621, 32'sd938, 32'sd1473, 32'sd907, 32'sd1390,
32'sd1398, 32'sd1712, 32'sd475, 32'sd1671, 32'sd659, 32'sd1301,
32'sd1417, 32'sd1558, 32'sd1357, 32'sd405, 32'sd881, 32'sd444,
32'sd202, 32'sd558, 32'sd389, 32'sd1216, 32'sd1044, 32'sd1404,
32'sd278, 32'sd804, 32'sd781, 32'sd1121, 32'sd829, 32'sd1217,
32'sd1029, 32'sd860, 32'sd1506, 32'sd1519, 32'sd1208, 32'sd962,
32'sd577, 32'sd1599, 32'sd1268, 32'sd777, 32'sd1342, 32'sd641,
32'sd759, 32'sd651, 32'sd1245, 32'sd519, 32'sd1107, 32'sd601,
32'sd1099, 32'sd1027, 32'sd493, 32'sd1692, 32'sd836, 32'sd2000,
32'sd1339, 32'sd1098, 32'sd1621, 32'sd1715, 32'sd1068, 32'sd211,
32'sd950, 32'sd1483, 32'sd1791, 32'sd348, 32'sd888, 32'sd1300,
32'sd187, 32'sd486, 32'sd881, 32'sd211, 32'sd1267, 32'sd1090,
32'sd1184, 32'sd1777, 32'sd269, 32'sd707, 32'sd1707, 32'sd1985,
32'sd114, 32'sd888, 32'sd1231, 32'sd762, 32'sd1252, 32'sd431,
32'sd373, 32'sd325, 32'sd166, 32'sd959, 32'sd1862, 32'sd1165,
32'sd568, 32'sd855, 32'sd125, 32'sd1017, 32'sd1067, 32'sd459,
32'sd1290, 32'sd1625, 32'sd111, 32'sd1547, 32'sd1264, 32'sd1532,
32'sd680, 32'sd1946, 32'sd830, 32'sd1755, 32'sd1080, 32'sd405,
32'sd981, 32'sd1994, 32'sd430, 32'sd1657, 32'sd641, 32'sd509,
32'sd1385, 32'sd1734, 32'sd1070, 32'sd894, 32'sd375, 32'sd1621,
32'sd1892, 32'sd1137, 32'sd1045, 32'sd432, 32'sd1164, 32'sd1348,
32'sd1971, 32'sd1049, 32'sd1297, 32'sd1751, 32'sd1060, 32'sd1361,
32'sd1314, 32'sd1107, 32'sd362, 32'sd276, 32'sd750, 32'sd984,
32'sd1206, 32'sd1516, 32'sd846, 32'sd1492, 32'sd1420, 32'sd682,
32'sd884, 32'sd1107, 32'sd1831, 32'sd1286, 32'sd948, 32'sd1605,
32'sd1576, 32'sd1663, 32'sd1930, 32'sd1096, 32'sd182, 32'sd1140,
32'sd1042, 32'sd1629, 32'sd1786, 32'sd898, 32'sd218, 32'sd1676,
32'sd1446, 32'sd1923, 32'sd1953, 32'sd1358, 32'sd1520, 32'sd591,
32'sd393, 32'sd1094, 32'sd1793, 32'sd746, 32'sd1128, 32'sd764,
32'sd292, 32'sd106, 32'sd710, 32'sd273, 32'sd1689, 32'sd1356,
32'sd1601, 32'sd1629, 32'sd1414, 32'sd488, 32'sd223, 32'sd225,
32'sd1395, 32'sd1892, 32'sd626, 32'sd1672, 32'sd1867, 32'sd1305,
32'sd1070, 32'sd1844, 32'sd1632, 32'sd714, 32'sd541, 32'sd1519,
32'sd271, 32'sd1151, 32'sd846, 32'sd1356, 32'sd453, 32'sd1149,
32'sd991, 32'sd1278, 32'sd1369, 32'sd230, 32'sd1359, 32'sd1911,
32'sd1798, 32'sd897, 32'sd553, 32'sd1353, 32'sd427, 32'sd1249,
32'sd495, 32'sd168, 32'sd1004, 32'sd978, 32'sd1627, 32'sd279,
32'sd1027, 32'sd1250, 32'sd1649, 32'sd786, 32'sd1642, 32'sd657,
32'sd793, 32'sd1498, 32'sd257, 32'sd484, 32'sd530, 32'sd1772,
32'sd1845, 32'sd263, 32'sd1250, 32'sd1607, 32'sd562, 32'sd1645,
32'sd375, 32'sd1003, 32'sd827, 32'sd359, 32'sd1682, 32'sd1601,
32'sd1230, 32'sd1430, 32'sd164, 32'sd1779, 32'sd1276, 32'sd297,
32'sd282, 32'sd1929, 32'sd1081, 32'sd1545, 32'sd1385, 32'sd1680,
32'sd554, 32'sd1168, 32'sd1080, 32'sd1055, 32'sd878, 32'sd451,
32'sd1935, 32'sd1109, 32'sd1556, 32'sd1554, 32'sd834, 32'sd1536,
32'sd480, 32'sd1539, 32'sd961, 32'sd865, 32'sd1770, 32'sd424,
32'sd1345, 32'sd1246, 32'sd880, 32'sd1071, 32'sd487, 32'sd1281,
32'sd1725, 32'sd1741, 32'sd997, 32'sd1965, 32'sd1611, 32'sd465,
32'sd884, 32'sd285, 32'sd325, 32'sd124, 32'sd339, 32'sd425,
32'sd1813, 32'sd1916, 32'sd1547, 32'sd1290, 32'sd1058, 32'sd1250,
32'sd186, 32'sd215, 32'sd1230, 32'sd1007, 32'sd321, 32'sd1020,
32'sd788, 32'sd1689, 32'sd451, 32'sd808, 32'sd1384, 32'sd1628,
32'sd709, 32'sd1723, 32'sd1924, 32'sd1027, 32'sd1267, 32'sd1619,
32'sd1098, 32'sd863, 32'sd1330, 32'sd1403, 32'sd660, 32'sd1863,
32'sd929, 32'sd543, 32'sd380, 32'sd1113, 32'sd644, 32'sd1045,
32'sd330, 32'sd1194, 32'sd207, 32'sd1147, 32'sd1821, 32'sd588,
32'sd1145, 32'sd305, 32'sd1576, 32'sd437, 32'sd1635, 32'sd962,
32'sd154, 32'sd744, 32'sd796, 32'sd1112, 32'sd1326, 32'sd1340,
32'sd784, 32'sd127, 32'sd1313, 32'sd1834, 32'sd321, 32'sd1974,
32'sd1844, 32'sd329, 32'sd1330, 32'sd1230, 32'sd749, 32'sd1048,
32'sd598, 32'sd772, 32'sd156, 32'sd1289, 32'sd1181, 32'sd1640,
32'sd335, 32'sd1900, 32'sd1371, 32'sd1153, 32'sd451, 32'sd1889,
32'sd960, 32'sd974, 32'sd778, 32'sd1962, 32'sd1150, 32'sd305,
32'sd792, 32'sd1339, 32'sd345, 32'sd1207, 32'sd1441, 32'sd1597,
32'sd768, 32'sd423, 32'sd1484, 32'sd934, 32'sd1791, 32'sd1211,
32'sd1484, 32'sd1603, 32'sd933, 32'sd1648, 32'sd470, 32'sd1786,
32'sd471, 32'sd1768, 32'sd154, 32'sd379, 32'sd170, 32'sd435,
32'sd327, 32'sd534, 32'sd1735, 32'sd236, 32'sd1987, 32'sd901,
32'sd1989, 32'sd223, 32'sd1224, 32'sd1118, 32'sd600, 32'sd1849,
32'sd1871, 32'sd815, 32'sd469, 32'sd506, 32'sd1351, 32'sd978,
32'sd656, 32'sd664, 32'sd1972, 32'sd1377, 32'sd1409, 32'sd1924,
32'sd1711, 32'sd1761, 32'sd240, 32'sd1592, 32'sd1350, 32'sd1784,
32'sd1137, 32'sd306, 32'sd1771, 32'sd1385, 32'sd1501, 32'sd861,
32'sd1810, 32'sd240, 32'sd946, 32'sd1342, 32'sd760, 32'sd433,
32'sd156, 32'sd179, 32'sd1538, 32'sd1826, 32'sd1356, 32'sd400,
32'sd1771, 32'sd576, 32'sd1668, 32'sd960, 32'sd1385, 32'sd1785,
32'sd744, 32'sd953, 32'sd1383, 32'sd1052, 32'sd681, 32'sd664,
32'sd1982, 32'sd1838, 32'sd596, 32'sd1234, 32'sd1114, 32'sd1679,
32'sd368, 32'sd613, 32'sd599, 32'sd1834, 32'sd1856, 32'sd1846,
32'sd672, 32'sd1572, 32'sd219, 32'sd1407, 32'sd1120, 32'sd1700,
32'sd975, 32'sd298, 32'sd420, 32'sd251, 32'sd1930, 32'sd794,
32'sd1146, 32'sd801, 32'sd1776, 32'sd1132, 32'sd418, 32'sd777,
32'sd1408, 32'sd1236, 32'sd539, 32'sd676, 32'sd213, 32'sd1824,
32'sd1215, 32'sd538, 32'sd1836, 32'sd1824, 32'sd122, 32'sd700,
32'sd504, 32'sd1535, 32'sd1054, 32'sd1037, 32'sd543, 32'sd1927,
32'sd1249, 32'sd348, 32'sd1041, 32'sd1791, 32'sd1670, 32'sd1238,
32'sd1517, 32'sd359, 32'sd502, 32'sd1066, 32'sd1075, 32'sd972,
32'sd1771, 32'sd659, 32'sd859, 32'sd133, 32'sd1550, 32'sd806,
32'sd1318, 32'sd1868, 32'sd150, 32'sd1052, 32'sd882, 32'sd1702,
32'sd1799, 32'sd1476, 32'sd541, 32'sd224, 32'sd233, 32'sd361,
32'sd835, 32'sd1928, 32'sd451, 32'sd1570, 32'sd1282, 32'sd734,
32'sd613, 32'sd484, 32'sd440, 32'sd217, 32'sd219, 32'sd1554,
32'sd345, 32'sd984, 32'sd1345, 32'sd1298, 32'sd454, 32'sd1563,
32'sd939, 32'sd1311, 32'sd162, 32'sd745, 32'sd538, 32'sd1207,
32'sd1837, 32'sd813, 32'sd695, 32'sd1407, 32'sd955, 32'sd1732,
32'sd1947, 32'sd875, 32'sd1891, 32'sd1189, 32'sd917, 32'sd1000,
32'sd768, 32'sd1030, 32'sd1708, 32'sd116, 32'sd232, 32'sd363,
32'sd337, 32'sd1843, 32'sd1250, 32'sd1347, 32'sd1384, 32'sd1181,
32'sd1878, 32'sd1575, 32'sd1756, 32'sd383, 32'sd892, 32'sd975,
32'sd409, 32'sd1494, 32'sd1085, 32'sd1642, 32'sd1784, 32'sd1603,
32'sd988, 32'sd1675, 32'sd856, 32'sd1659, 32'sd1763, 32'sd1933,
32'sd837, 32'sd999, 32'sd901, 32'sd1542, 32'sd319, 32'sd1893,
32'sd1856, 32'sd1177, 32'sd700, 32'sd466, 32'sd1905, 32'sd872,
32'sd850, 32'sd953, 32'sd800, 32'sd982, 32'sd750, 32'sd191,
32'sd148, 32'sd1332, 32'sd1697, 32'sd881, 32'sd1820, 32'sd578,
32'sd156, 32'sd760, 32'sd1177, 32'sd1075, 32'sd1019, 32'sd402,
32'sd790, 32'sd427, 32'sd1802, 32'sd1107, 32'sd353, 32'sd1620,
32'sd1857, 32'sd1519, 32'sd545, 32'sd772, 32'sd612, 32'sd953,
32'sd767, 32'sd1454, 32'sd296, 32'sd420, 32'sd1232, 32'sd1126,
32'sd1139, 32'sd932, 32'sd971, 32'sd1060, 32'sd378, 32'sd1788,
32'sd120, 32'sd274, 32'sd870, 32'sd799, 32'sd443, 32'sd1356,
32'sd1151, 32'sd1436, 32'sd127, 32'sd1493, 32'sd670, 32'sd656,
32'sd105, 32'sd1172, 32'sd776, 32'sd1619, 32'sd1845, 32'sd403,
32'sd1121, 32'sd1412, 32'sd1074, 32'sd1416, 32'sd1274, 32'sd1943,
32'sd536, 32'sd286, 32'sd256, 32'sd526, 32'sd1042, 32'sd1725,
32'sd1951, 32'sd142, 32'sd1165, 32'sd759, 32'sd1808, 32'sd744,
32'sd1496, 32'sd1167, 32'sd425, 32'sd1516, 32'sd1433, 32'sd341,
32'sd627, 32'sd248, 32'sd525, 32'sd487, 32'sd119, 32'sd1665,
32'sd440, 32'sd1546, 32'sd1551, 32'sd237, 32'sd1112, 32'sd1625,
32'sd913, 32'sd1107, 32'sd1321, 32'sd1531, 32'sd1022, 32'sd1034,
32'sd218, 32'sd1951, 32'sd993, 32'sd690, 32'sd1254, 32'sd973,
32'sd1364, 32'sd1675, 32'sd1914, 32'sd1666, 32'sd1893, 32'sd170,
32'sd493, 32'sd414, 32'sd909, 32'sd1630, 32'sd1616, 32'sd385,
32'sd373, 32'sd676, 32'sd1327, 32'sd1721, 32'sd1337, 32'sd407,
32'sd952, 32'sd544, 32'sd1166, 32'sd1771, 32'sd1757, 32'sd1564,
32'sd1225, 32'sd1173, 32'sd693, 32'sd1728, 32'sd297, 32'sd1858,
32'sd579, 32'sd1991, 32'sd314, 32'sd1158, 32'sd1517, 32'sd1535,
32'sd1957, 32'sd569, 32'sd1447, 32'sd1295, 32'sd611, 32'sd1727,
32'sd952, 32'sd800, 32'sd1220, 32'sd765, 32'sd1677, 32'sd683,
32'sd1646, 32'sd123, 32'sd1114, 32'sd1438, 32'sd1750, 32'sd1697,
32'sd1139, 32'sd1506, 32'sd1890, 32'sd1052, 32'sd1460, 32'sd1111,
32'sd1595, 32'sd1933, 32'sd1103, 32'sd666, 32'sd1732, 32'sd1497,
32'sd377, 32'sd1389, 32'sd120, 32'sd867, 32'sd443, 32'sd148,
32'sd1993, 32'sd706, 32'sd1382, 32'sd1298, 32'sd223, 32'sd1873,
32'sd1790, 32'sd623, 32'sd870, 32'sd861, 32'sd688, 32'sd970,
32'sd1425, 32'sd1100, 32'sd863, 32'sd626, 32'sd771, 32'sd1733,
32'sd1045, 32'sd1455, 32'sd1166, 32'sd1520, 32'sd783, 32'sd980,
32'sd1162, 32'sd1619, 32'sd918, 32'sd401, 32'sd1683, 32'sd1115,
32'sd656, 32'sd1303, 32'sd1822, 32'sd355, 32'sd313, 32'sd1371,
32'sd883, 32'sd1822, 32'sd919, 32'sd1297, 32'sd1521, 32'sd744,
32'sd1080, 32'sd972, 32'sd1500, 32'sd1731, 32'sd1228, 32'sd144,
32'sd1521, 32'sd1281, 32'sd489, 32'sd509, 32'sd1375, 32'sd1124,
32'sd699, 32'sd821, 32'sd1532, 32'sd1174, 32'sd810, 32'sd1942,
32'sd1599, 32'sd602, 32'sd597, 32'sd1673, 32'sd145, 32'sd1939,
32'sd886, 32'sd973, 32'sd900, 32'sd141, 32'sd1053, 32'sd1595,
32'sd662, 32'sd1393, 32'sd126, 32'sd1761, 32'sd311, 32'sd1395,
32'sd1659, 32'sd434, 32'sd1353, 32'sd1031, 32'sd126, 32'sd447,
32'sd1593, 32'sd1737, 32'sd350, 32'sd1513, 32'sd1566, 32'sd919,
32'sd1432, 32'sd1113, 32'sd1800, 32'sd133, 32'sd157, 32'sd718,
32'sd974, 32'sd534, 32'sd975, 32'sd871, 32'sd346, 32'sd1081,
32'sd1487, 32'sd948, 32'sd1536, 32'sd242, 32'sd1398, 32'sd475,
32'sd1667, 32'sd1647, 32'sd799, 32'sd581, 32'sd1897, 32'sd1425,
32'sd772, 32'sd1368, 32'sd1378, 32'sd1292, 32'sd1727, 32'sd886,
32'sd943, 32'sd984, 32'sd795, 32'sd824, 32'sd555, 32'sd447,
32'sd1839, 32'sd1782, 32'sd1404, 32'sd847, 32'sd1160, 32'sd1811,
32'sd418, 32'sd1712, 32'sd1627, 32'sd1871, 32'sd303, 32'sd711,
32'sd1365, 32'sd475, 32'sd702, 32'sd577, 32'sd1836, 32'sd606,
32'sd1816, 32'sd1022, 32'sd295, 32'sd692, 32'sd1437, 32'sd1381,
32'sd1763, 32'sd1577, 32'sd1074, 32'sd1938, 32'sd1512, 32'sd1952,
32'sd201, 32'sd1368, 32'sd381, 32'sd257, 32'sd1207, 32'sd1520,
32'sd1771, 32'sd402, 32'sd387, 32'sd956, 32'sd361, 32'sd200,
32'sd364, 32'sd327, 32'sd314, 32'sd916, 32'sd1614, 32'sd886,
32'sd1841, 32'sd1286, 32'sd486, 32'sd1561, 32'sd1027, 32'sd1156,
32'sd1423, 32'sd1217, 32'sd1099, 32'sd1847, 32'sd1475, 32'sd1429,
32'sd1738, 32'sd250, 32'sd1743, 32'sd1680, 32'sd891, 32'sd355,
32'sd190, 32'sd1578, 32'sd208, 32'sd792, 32'sd993, 32'sd1877,
32'sd1784, 32'sd1752, 32'sd1802, 32'sd802, 32'sd1961, 32'sd725,
32'sd1011, 32'sd272, 32'sd651, 32'sd156, 32'sd216, 32'sd102,
32'sd1069, 32'sd1549, 32'sd1533, 32'sd1842, 32'sd1056, 32'sd522,
32'sd806, 32'sd1898, 32'sd727, 32'sd1621, 32'sd1982, 32'sd1273,
32'sd676, 32'sd1521, 32'sd1598, 32'sd995, 32'sd498, 32'sd1855,
32'sd618, 32'sd685, 32'sd1858, 32'sd341, 32'sd129, 32'sd1415,
32'sd1748, 32'sd623, 32'sd1477, 32'sd506, 32'sd209, 32'sd1085,
32'sd1346, 32'sd1122, 32'sd1685, 32'sd1609, 32'sd1517, 32'sd1503,
32'sd857, 32'sd798, 32'sd437, 32'sd521, 32'sd1991, 32'sd1877,
32'sd684, 32'sd1846, 32'sd1884, 32'sd1591, 32'sd1081, 32'sd1691,
32'sd853, 32'sd1263, 32'sd1632, 32'sd914, 32'sd681, 32'sd1727,
32'sd1170, 32'sd906, 32'sd578, 32'sd193, 32'sd1376, 32'sd753,
32'sd983, 32'sd731, 32'sd1856, 32'sd936, 32'sd177, 32'sd1483,
32'sd167, 32'sd1472, 32'sd1111, 32'sd1856, 32'sd780, 32'sd1529,
32'sd504, 32'sd1783, 32'sd141, 32'sd1963, 32'sd541, 32'sd1187,
32'sd1311, 32'sd547, 32'sd1276, 32'sd680, 32'sd1449, 32'sd587,
32'sd1182, 32'sd1280, 32'sd1769, 32'sd243, 32'sd1220, 32'sd721,
32'sd496, 32'sd1049, 32'sd454, 32'sd1871, 32'sd828, 32'sd731,
32'sd876, 32'sd858, 32'sd1009, 32'sd1546, 32'sd468, 32'sd254,
32'sd681, 32'sd237, 32'sd549, 32'sd722, 32'sd804, 32'sd1532,
32'sd680, 32'sd949, 32'sd496, 32'sd1128, 32'sd946, 32'sd1677,
32'sd1603, 32'sd878, 32'sd159, 32'sd625, 32'sd279, 32'sd1796,
32'sd1161, 32'sd488, 32'sd1938, 32'sd568, 32'sd412, 32'sd1882,
32'sd120, 32'sd1693, 32'sd1522, 32'sd203, 32'sd573, 32'sd1181,
32'sd1359, 32'sd1300, 32'sd1142, 32'sd376, 32'sd758, 32'sd1315,
32'sd1812, 32'sd805, 32'sd216, 32'sd685, 32'sd1955, 32'sd918,
32'sd1512, 32'sd510, 32'sd133, 32'sd373, 32'sd1778, 32'sd1888,
32'sd340, 32'sd1562, 32'sd1400, 32'sd1443, 32'sd965, 32'sd1877,
32'sd1843, 32'sd120, 32'sd630, 32'sd851, 32'sd1810, 32'sd410,
32'sd657, 32'sd1135, 32'sd1752, 32'sd301, 32'sd1624, 32'sd1739,
32'sd1649, 32'sd1286, 32'sd1592, 32'sd478, 32'sd1168, 32'sd1160,
32'sd1119, 32'sd189, 32'sd1212, 32'sd1315, 32'sd1653, 32'sd495,
32'sd1471, 32'sd1013, 32'sd834, 32'sd419, 32'sd1128, 32'sd1518,
32'sd1318, 32'sd967, 32'sd629, 32'sd1025, 32'sd237, 32'sd365,
32'sd1342, 32'sd1767, 32'sd644, 32'sd960, 32'sd475, 32'sd770,
32'sd1693, 32'sd712, 32'sd342, 32'sd603, 32'sd1415, 32'sd1578,
32'sd847, 32'sd1582, 32'sd662, 32'sd1635, 32'sd212, 32'sd191,
32'sd705, 32'sd1189, 32'sd308, 32'sd914, 32'sd1563, 32'sd529,
32'sd1135, 32'sd1008, 32'sd1580, 32'sd321, 32'sd163, 32'sd834,
32'sd1503, 32'sd1100, 32'sd497, 32'sd536, 32'sd804, 32'sd1195,
32'sd441, 32'sd183, 32'sd1427, 32'sd364, 32'sd236, 32'sd1839,
32'sd944, 32'sd922, 32'sd1727, 32'sd918, 32'sd695, 32'sd1637,
32'sd926, 32'sd891, 32'sd1209, 32'sd1595, 32'sd765, 32'sd805,
32'sd451, 32'sd187, 32'sd1544, 32'sd1512, 32'sd1117, 32'sd156,
32'sd1181, 32'sd233, 32'sd1895, 32'sd626, 32'sd867, 32'sd1667,
32'sd1533, 32'sd1395, 32'sd437, 32'sd1516, 32'sd1989, 32'sd1631,
32'sd1588, 32'sd1628, 32'sd1288, 32'sd1738, 32'sd235, 32'sd1208,
32'sd1948, 32'sd1114, 32'sd435, 32'sd310, 32'sd590, 32'sd426,
32'sd1342, 32'sd1723, 32'sd1206, 32'sd1865, 32'sd345, 32'sd1708,
32'sd350, 32'sd175, 32'sd1877, 32'sd649, 32'sd1282, 32'sd376,
32'sd563, 32'sd889, 32'sd1317, 32'sd721, 32'sd1326, 32'sd356,
32'sd289, 32'sd1787, 32'sd964, 32'sd249, 32'sd1801, 32'sd192,
32'sd1756, 32'sd1176, 32'sd1878, 32'sd1830, 32'sd1526, 32'sd1688,
32'sd749, 32'sd1100, 32'sd1708, 32'sd1787, 32'sd638, 32'sd727,
32'sd1384, 32'sd1039, 32'sd517, 32'sd1971, 32'sd1729, 32'sd103,
32'sd1274, 32'sd323, 32'sd639, 32'sd1950, 32'sd1446, 32'sd1359,
32'sd936, 32'sd269, 32'sd549, 32'sd1613, 32'sd1717, 32'sd1510,
32'sd1888, 32'sd599, 32'sd473, 32'sd686, 32'sd332, 32'sd432,
32'sd1146, 32'sd1241, 32'sd578, 32'sd1177, 32'sd1800, 32'sd1936,
32'sd1754, 32'sd1665, 32'sd207, 32'sd294, 32'sd1392, 32'sd1090,
32'sd1118, 32'sd867, 32'sd1079, 32'sd1370, 32'sd807, 32'sd1671,
32'sd491, 32'sd794, 32'sd859, 32'sd1693, 32'sd1745, 32'sd1384,
32'sd102, 32'sd1511, 32'sd1723, 32'sd810, 32'sd351, 32'sd1503,
32'sd1007, 32'sd1155, 32'sd1431, 32'sd222, 32'sd622, 32'sd779,
32'sd1328, 32'sd974, 32'sd423, 32'sd314, 32'sd1101, 32'sd643,
32'sd1217, 32'sd360, 32'sd1309, 32'sd480, 32'sd1332, 32'sd424,
32'sd443, 32'sd1754, 32'sd1329, 32'sd1174, 32'sd824, 32'sd1932,
32'sd578, 32'sd148, 32'sd1533, 32'sd1890, 32'sd730, 32'sd1844,
32'sd1763, 32'sd770, 32'sd1758, 32'sd1664, 32'sd424, 32'sd133,
32'sd704, 32'sd192, 32'sd1694, 32'sd827, 32'sd398, 32'sd1564,
32'sd402, 32'sd1374, 32'sd905, 32'sd257, 32'sd1979, 32'sd1477,
32'sd1648, 32'sd1857, 32'sd1315, 32'sd485, 32'sd102, 32'sd898,
32'sd339, 32'sd335, 32'sd309, 32'sd1511, 32'sd245, 32'sd312,
32'sd1955, 32'sd704, 32'sd1562, 32'sd1112, 32'sd1183, 32'sd587,
32'sd1045, 32'sd1826, 32'sd710, 32'sd1809, 32'sd675, 32'sd772,
32'sd615, 32'sd1578, 32'sd1552, 32'sd785, 32'sd542, 32'sd706,
32'sd1844, 32'sd204, 32'sd368, 32'sd612, 32'sd616, 32'sd1138,
32'sd605, 32'sd1970, 32'sd1626, 32'sd846, 32'sd1214, 32'sd1925,
32'sd1494, 32'sd604, 32'sd1925, 32'sd1411, 32'sd138, 32'sd670,
32'sd1922, 32'sd1788, 32'sd1440, 32'sd1472, 32'sd1482, 32'sd1743,
32'sd1877, 32'sd224, 32'sd1052, 32'sd1723, 32'sd428, 32'sd509,
32'sd1676, 32'sd1420, 32'sd804, 32'sd1461, 32'sd1029, 32'sd1309,
32'sd1089, 32'sd1893, 32'sd1029, 32'sd271, 32'sd1842, 32'sd1092,
32'sd114, 32'sd1183, 32'sd146, 32'sd518, 32'sd1116, 32'sd958,
32'sd946, 32'sd1000, 32'sd908, 32'sd1924, 32'sd472, 32'sd1504,
32'sd420, 32'sd662, 32'sd1644, 32'sd1138, 32'sd690, 32'sd1820,
32'sd851, 32'sd964, 32'sd1146, 32'sd430, 32'sd1486, 32'sd1234,
32'sd885, 32'sd469, 32'sd1664, 32'sd780, 32'sd1880, 32'sd1704,
32'sd584, 32'sd150, 32'sd602, 32'sd219, 32'sd1662, 32'sd1664,
32'sd1214, 32'sd1185, 32'sd841, 32'sd1053, 32'sd354, 32'sd1248,
32'sd371, 32'sd1408, 32'sd318, 32'sd1230, 32'sd1629, 32'sd701,
32'sd1084, 32'sd1656, 32'sd747, 32'sd1560, 32'sd382, 32'sd671,
32'sd1271, 32'sd1339, 32'sd969, 32'sd682, 32'sd1756, 32'sd148,
32'sd154, 32'sd931, 32'sd875, 32'sd1022, 32'sd1689, 32'sd1828,
32'sd1211, 32'sd1846, 32'sd1708, 32'sd982, 32'sd1582, 32'sd1233,
32'sd1549, 32'sd1665, 32'sd691, 32'sd1229, 32'sd1080, 32'sd308,
32'sd460, 32'sd1166, 32'sd670, 32'sd680, 32'sd1741, 32'sd1592,
32'sd751, 32'sd1692, 32'sd828, 32'sd1273, 32'sd1834, 32'sd1036,
32'sd1432, 32'sd1111, 32'sd226, 32'sd1239, 32'sd271, 32'sd1300,
32'sd438, 32'sd1139, 32'sd1761, 32'sd1067, 32'sd1282, 32'sd249,
32'sd1808, 32'sd1720, 32'sd995, 32'sd1888, 32'sd1000, 32'sd1344,
32'sd723, 32'sd775, 32'sd1101, 32'sd1871, 32'sd812, 32'sd589,
32'sd304, 32'sd868, 32'sd1321, 32'sd262, 32'sd1470, 32'sd691,
32'sd757, 32'sd694, 32'sd157, 32'sd1568, 32'sd1703, 32'sd904,
32'sd1270, 32'sd1494, 32'sd1365, 32'sd1237, 32'sd1459, 32'sd466,
32'sd232, 32'sd149, 32'sd627, 32'sd1598, 32'sd623, 32'sd1680,
32'sd737, 32'sd1141, 32'sd1709, 32'sd317, 32'sd709, 32'sd1193,
32'sd564, 32'sd1116, 32'sd487, 32'sd484, 32'sd1427, 32'sd617,
32'sd137, 32'sd1465, 32'sd599, 32'sd1016, 32'sd1443, 32'sd412,
32'sd1017, 32'sd958, 32'sd707, 32'sd1254, 32'sd646, 32'sd198,
32'sd1019, 32'sd730, 32'sd1846, 32'sd429, 32'sd1481, 32'sd1671,
32'sd728, 32'sd1950, 32'sd722, 32'sd539, 32'sd365, 32'sd1398,
32'sd1823, 32'sd1799, 32'sd227, 32'sd895, 32'sd1231, 32'sd1273,
32'sd1450, 32'sd1243, 32'sd569, 32'sd1092, 32'sd1480, 32'sd1901,
32'sd1523, 32'sd766, 32'sd1346, 32'sd310, 32'sd1394, 32'sd689,
32'sd1469, 32'sd318, 32'sd1967, 32'sd801, 32'sd1379, 32'sd874,
32'sd1237, 32'sd1747, 32'sd1249, 32'sd1802, 32'sd1441, 32'sd1689,
32'sd808, 32'sd1534, 32'sd1431, 32'sd1979, 32'sd1076, 32'sd1590,
32'sd1696, 32'sd879, 32'sd1803, 32'sd575, 32'sd178, 32'sd733,
32'sd1107, 32'sd571, 32'sd1068, 32'sd380, 32'sd161, 32'sd1495,
32'sd928, 32'sd394, 32'sd1416, 32'sd943, 32'sd1090, 32'sd455,
32'sd170, 32'sd1942, 32'sd334, 32'sd1953, 32'sd317, 32'sd1035,
32'sd731, 32'sd248, 32'sd387, 32'sd807, 32'sd1347, 32'sd551,
32'sd1176, 32'sd339, 32'sd646, 32'sd1843, 32'sd133, 32'sd151,
32'sd1143, 32'sd369, 32'sd776, 32'sd1316, 32'sd1454, 32'sd1615,
32'sd1747, 32'sd1977, 32'sd842, 32'sd897, 32'sd323, 32'sd694,
32'sd1776, 32'sd1139, 32'sd1418, 32'sd150, 32'sd786, 32'sd1301,
32'sd1409, 32'sd460, 32'sd1715, 32'sd1727, 32'sd651, 32'sd1291,
32'sd1261, 32'sd1489, 32'sd302, 32'sd1782, 32'sd726, 32'sd1219,
32'sd1033, 32'sd1430, 32'sd1615, 32'sd340, 32'sd1294, 32'sd1052,
32'sd1387, 32'sd159, 32'sd313, 32'sd702, 32'sd1067, 32'sd1623,
32'sd1055, 32'sd1896, 32'sd1917, 32'sd297, 32'sd1804, 32'sd675,
32'sd1044, 32'sd1753, 32'sd1241, 32'sd1968, 32'sd507, 32'sd1770,
32'sd1508, 32'sd1860, 32'sd1034, 32'sd1796, 32'sd914, 32'sd1116,
32'sd1801, 32'sd1901, 32'sd1177, 32'sd484, 32'sd162, 32'sd947,
32'sd378, 32'sd1433, 32'sd1157, 32'sd689, 32'sd611, 32'sd709,
32'sd1045, 32'sd782, 32'sd1646, 32'sd1037, 32'sd1168, 32'sd1735,
32'sd117, 32'sd1755, 32'sd1618, 32'sd1073, 32'sd1823, 32'sd737,
32'sd537, 32'sd418, 32'sd443, 32'sd1901, 32'sd329, 32'sd318,
32'sd346, 32'sd1675, 32'sd1245, 32'sd1910, 32'sd1372, 32'sd1625,
32'sd584, 32'sd134, 32'sd1688, 32'sd1541, 32'sd825, 32'sd1418,
32'sd313, 32'sd327, 32'sd542, 32'sd1417, 32'sd351, 32'sd550,
32'sd1017, 32'sd362, 32'sd1792, 32'sd731, 32'sd802, 32'sd1013,
32'sd212, 32'sd1960, 32'sd1835, 32'sd362, 32'sd158, 32'sd1823,
32'sd1899, 32'sd363, 32'sd1270, 32'sd1596, 32'sd1909, 32'sd1036,
32'sd402, 32'sd145, 32'sd1264, 32'sd605, 32'sd191, 32'sd519,
32'sd387, 32'sd663, 32'sd1176, 32'sd999, 32'sd1857, 32'sd1569,
32'sd946, 32'sd703, 32'sd1341, 32'sd1500, 32'sd1317, 32'sd1470,
32'sd361, 32'sd1944, 32'sd368, 32'sd1539, 32'sd625, 32'sd290,
32'sd578, 32'sd1225, 32'sd374, 32'sd1375, 32'sd166, 32'sd1308,
32'sd1252, 32'sd1714, 32'sd587, 32'sd776, 32'sd738, 32'sd1629,
32'sd172, 32'sd978, 32'sd1215, 32'sd226, 32'sd1377, 32'sd1742,
32'sd869, 32'sd1834, 32'sd1062, 32'sd1325, 32'sd924, 32'sd1659,
32'sd241, 32'sd227, 32'sd1183, 32'sd866, 32'sd1953, 32'sd1822,
32'sd354, 32'sd1855, 32'sd1442, 32'sd405, 32'sd1883, 32'sd643,
32'sd1645, 32'sd549, 32'sd1212, 32'sd1226, 32'sd968, 32'sd1173,
32'sd910, 32'sd536, 32'sd362, 32'sd1555, 32'sd1369, 32'sd1684,
32'sd1436, 32'sd590, 32'sd1285, 32'sd834, 32'sd701, 32'sd1069,
32'sd231, 32'sd1497, 32'sd1323, 32'sd1586, 32'sd1281, 32'sd1542,
32'sd1565, 32'sd1043, 32'sd1944, 32'sd986, 32'sd386, 32'sd981,
32'sd334, 32'sd1620, 32'sd942, 32'sd1010, 32'sd145, 32'sd773,
32'sd1113, 32'sd240, 32'sd1493, 32'sd211, 32'sd991, 32'sd1562,
32'sd1518, 32'sd1870, 32'sd1097, 32'sd1118, 32'sd583, 32'sd364,
32'sd1164, 32'sd1730, 32'sd471, 32'sd1837, 32'sd1682, 32'sd1282,
32'sd1213, 32'sd1252, 32'sd1323, 32'sd457, 32'sd1321, 32'sd759,
32'sd983, 32'sd1833, 32'sd882, 32'sd556, 32'sd724, 32'sd1155,
32'sd194, 32'sd586, 32'sd1398, 32'sd175, 32'sd951, 32'sd1580,
32'sd1764, 32'sd1450, 32'sd1705, 32'sd1401, 32'sd1365, 32'sd1818,
32'sd401, 32'sd1177, 32'sd1152, 32'sd558, 32'sd329, 32'sd1410,
32'sd1479, 32'sd902, 32'sd1070, 32'sd669, 32'sd1823, 32'sd1478,
32'sd699, 32'sd1243, 32'sd585, 32'sd622, 32'sd1796, 32'sd1418,
32'sd836, 32'sd640, 32'sd652, 32'sd812, 32'sd1462, 32'sd643,
32'sd661, 32'sd729, 32'sd1372, 32'sd481, 32'sd1162, 32'sd559,
32'sd1586, 32'sd1262, 32'sd269, 32'sd201, 32'sd1811, 32'sd1125,
32'sd457, 32'sd327, 32'sd992, 32'sd1845, 32'sd235, 32'sd1957,
32'sd229, 32'sd1370, 32'sd1726, 32'sd1413, 32'sd1147, 32'sd1417,
32'sd488, 32'sd236, 32'sd112, 32'sd456, 32'sd1081, 32'sd1819,
32'sd576, 32'sd1612, 32'sd1888, 32'sd1205, 32'sd1219, 32'sd277,
32'sd254, 32'sd408, 32'sd1692, 32'sd681, 32'sd628, 32'sd1175,
32'sd112, 32'sd1865, 32'sd911, 32'sd372, 32'sd1539, 32'sd1380,
32'sd691, 32'sd1177, 32'sd305, 32'sd123, 32'sd254, 32'sd263,
32'sd1117, 32'sd1630, 32'sd1743, 32'sd1835, 32'sd1019, 32'sd1794,
32'sd1909, 32'sd930, 32'sd1126, 32'sd1996, 32'sd1913, 32'sd874,
32'sd1365, 32'sd536, 32'sd595, 32'sd1581, 32'sd243, 32'sd403,
32'sd1539, 32'sd1323, 32'sd1892, 32'sd1501, 32'sd524, 32'sd1543,
32'sd1721, 32'sd1495, 32'sd938, 32'sd787, 32'sd1524, 32'sd1464,
32'sd1831, 32'sd134, 32'sd1339, 32'sd246, 32'sd1265, 32'sd602,
32'sd124, 32'sd1708, 32'sd661, 32'sd1041, 32'sd759, 32'sd1823,
32'sd966, 32'sd973, 32'sd143, 32'sd863, 32'sd1835, 32'sd777,
32'sd1637, 32'sd736, 32'sd1821, 32'sd661, 32'sd1033, 32'sd1645,
32'sd1461, 32'sd1420, 32'sd645, 32'sd221, 32'sd1747, 32'sd1961,
32'sd277, 32'sd1626, 32'sd845, 32'sd1147, 32'sd1976, 32'sd1513,
32'sd499, 32'sd1393, 32'sd1706, 32'sd381, 32'sd1818, 32'sd1620,
32'sd398, 32'sd1114, 32'sd1328, 32'sd1109, 32'sd1515, 32'sd953,
32'sd381, 32'sd221, 32'sd213, 32'sd1690, 32'sd1166, 32'sd1152,
32'sd1026, 32'sd445, 32'sd882, 32'sd284, 32'sd1496, 32'sd149,
32'sd1250, 32'sd1493, 32'sd483, 32'sd1353, 32'sd533, 32'sd274,
32'sd818, 32'sd1830, 32'sd1568, 32'sd221, 32'sd1340, 32'sd711,
32'sd1559, 32'sd586, 32'sd1690, 32'sd1109, 32'sd520, 32'sd1185,
32'sd691, 32'sd1365, 32'sd495, 32'sd265, 32'sd1022, 32'sd1635,
32'sd461, 32'sd1454, 32'sd1436, 32'sd1310, 32'sd664, 32'sd1583,
32'sd820, 32'sd230, 32'sd1654, 32'sd1072, 32'sd972, 32'sd1564,
32'sd1474, 32'sd1033, 32'sd1758, 32'sd389, 32'sd1434, 32'sd503,
32'sd1088, 32'sd100, 32'sd540, 32'sd491, 32'sd1149, 32'sd457,
32'sd440, 32'sd1540, 32'sd1930, 32'sd333, 32'sd1736, 32'sd668,
32'sd248, 32'sd1437, 32'sd1272, 32'sd1163, 32'sd1452, 32'sd1012,
32'sd271, 32'sd590, 32'sd751, 32'sd1460, 32'sd658, 32'sd1999,
32'sd196, 32'sd1776, 32'sd230, 32'sd389, 32'sd986, 32'sd327,
32'sd783, 32'sd917, 32'sd284, 32'sd139, 32'sd1681, 32'sd413,
32'sd1706, 32'sd1819, 32'sd1583, 32'sd1910, 32'sd1609, 32'sd852,
32'sd727, 32'sd1090, 32'sd1615, 32'sd974, 32'sd1003, 32'sd1156,
32'sd1366, 32'sd273, 32'sd1448, 32'sd423, 32'sd1683, 32'sd310,
32'sd1615, 32'sd1774, 32'sd671, 32'sd156, 32'sd489, 32'sd1832,
32'sd1263, 32'sd1111, 32'sd140, 32'sd1021, 32'sd1991, 32'sd1642,
32'sd1127, 32'sd1153, 32'sd376, 32'sd1456, 32'sd1184, 32'sd526,
32'sd582, 32'sd657, 32'sd449, 32'sd782, 32'sd1940, 32'sd1647,
32'sd849, 32'sd119, 32'sd1125, 32'sd1436, 32'sd1661, 32'sd1313,
32'sd468, 32'sd1599, 32'sd1605, 32'sd808, 32'sd794, 32'sd764,
32'sd1270, 32'sd1676, 32'sd811, 32'sd1310, 32'sd1874, 32'sd1830,
32'sd1976, 32'sd1700, 32'sd286, 32'sd877, 32'sd598, 32'sd1430,
32'sd742, 32'sd1920, 32'sd366, 32'sd464, 32'sd911, 32'sd1261,
32'sd1172, 32'sd708, 32'sd887, 32'sd892, 32'sd1102, 32'sd998,
32'sd380, 32'sd1219, 32'sd699, 32'sd1536, 32'sd254, 32'sd1548,
32'sd1398, 32'sd1667, 32'sd448, 32'sd1379, 32'sd512, 32'sd1009,
32'sd1759, 32'sd1272, 32'sd981, 32'sd596, 32'sd826, 32'sd1050,
32'sd743, 32'sd1790, 32'sd938, 32'sd852, 32'sd338, 32'sd1311,
32'sd871, 32'sd816, 32'sd898, 32'sd487, 32'sd711, 32'sd786,
32'sd1278, 32'sd610, 32'sd588, 32'sd341, 32'sd114, 32'sd208,
32'sd205, 32'sd687, 32'sd1042, 32'sd1897, 32'sd1036, 32'sd1009,
32'sd1452, 32'sd853, 32'sd852, 32'sd295, 32'sd711, 32'sd965,
32'sd440, 32'sd1570, 32'sd1085, 32'sd1890, 32'sd164, 32'sd1730,
32'sd1100, 32'sd1348, 32'sd1012, 32'sd1240, 32'sd950, 32'sd508,
32'sd1847, 32'sd1482, 32'sd1781, 32'sd252, 32'sd1807, 32'sd966,
32'sd655, 32'sd944, 32'sd1231, 32'sd1131, 32'sd1636, 32'sd698,
32'sd667, 32'sd1358, 32'sd1207, 32'sd828, 32'sd1723, 32'sd1025,
32'sd841, 32'sd1510, 32'sd1375, 32'sd1547, 32'sd1272, 32'sd1799,
32'sd1007, 32'sd1101, 32'sd364, 32'sd217, 32'sd1120, 32'sd1161,
32'sd1345, 32'sd363, 32'sd1292, 32'sd1958, 32'sd1149, 32'sd1289,
32'sd1152, 32'sd1299, 32'sd1680, 32'sd448, 32'sd227, 32'sd933,
32'sd191, 32'sd1735, 32'sd1095, 32'sd1865, 32'sd103, 32'sd948,
32'sd1544, 32'sd1426, 32'sd234, 32'sd1148, 32'sd662, 32'sd1360,
32'sd952, 32'sd854, 32'sd706, 32'sd959, 32'sd1126, 32'sd1074,
32'sd1554, 32'sd564, 32'sd1186, 32'sd868, 32'sd225, 32'sd956,
32'sd1659, 32'sd391, 32'sd138, 32'sd319, 32'sd1848, 32'sd1339,
32'sd636, 32'sd598, 32'sd714, 32'sd1317, 32'sd179, 32'sd895,
32'sd414, 32'sd1887, 32'sd1671, 32'sd1059, 32'sd801, 32'sd1566,
32'sd440, 32'sd795, 32'sd559, 32'sd1315, 32'sd1053, 32'sd170,
32'sd1821, 32'sd1638, 32'sd564, 32'sd913, 32'sd1950, 32'sd858,
32'sd1912, 32'sd931, 32'sd1893, 32'sd1841, 32'sd409, 32'sd821,
32'sd434, 32'sd429, 32'sd1096, 32'sd164, 32'sd1871, 32'sd597,
32'sd1625, 32'sd1895, 32'sd775, 32'sd202, 32'sd1005, 32'sd442,
32'sd723, 32'sd1361, 32'sd792, 32'sd1808, 32'sd1725, 32'sd1582,
32'sd1463, 32'sd101, 32'sd843, 32'sd1947, 32'sd1975, 32'sd1599,
32'sd1094, 32'sd1109, 32'sd1669, 32'sd773, 32'sd392, 32'sd1888,
32'sd171, 32'sd1938, 32'sd1839, 32'sd395, 32'sd1283, 32'sd1857,
32'sd1515, 32'sd978, 32'sd1489, 32'sd1726, 32'sd1689, 32'sd804,
32'sd615, 32'sd233, 32'sd303, 32'sd1439, 32'sd1765, 32'sd869,
32'sd1296, 32'sd1106, 32'sd582, 32'sd1592, 32'sd1314, 32'sd905,
32'sd1239, 32'sd555, 32'sd1399, 32'sd353, 32'sd925, 32'sd873,
32'sd198, 32'sd381, 32'sd435, 32'sd1164, 32'sd1934, 32'sd1243,
32'sd1726, 32'sd1836, 32'sd160, 32'sd789, 32'sd162, 32'sd489,
32'sd1350, 32'sd491, 32'sd1145, 32'sd1419, 32'sd1603, 32'sd269,
32'sd821, 32'sd125, 32'sd1992, 32'sd216, 32'sd558, 32'sd1572,
32'sd1280, 32'sd1377, 32'sd1699, 32'sd1243, 32'sd849, 32'sd492,
32'sd1997, 32'sd1507, 32'sd177, 32'sd155, 32'sd894, 32'sd406,
32'sd1283, 32'sd1144, 32'sd527, 32'sd1437, 32'sd1467, 32'sd153,
32'sd1380, 32'sd1969, 32'sd547, 32'sd1468, 32'sd545, 32'sd388,
32'sd1334, 32'sd731, 32'sd337, 32'sd1565, 32'sd1511, 32'sd1658,
32'sd896, 32'sd695, 32'sd567, 32'sd1271, 32'sd698, 32'sd815,
32'sd978, 32'sd133, 32'sd1667, 32'sd593, 32'sd1288, 32'sd314,
32'sd1108, 32'sd1682, 32'sd470, 32'sd1690, 32'sd139, 32'sd627,
32'sd296, 32'sd950, 32'sd391, 32'sd1090, 32'sd134, 32'sd652,
32'sd1750, 32'sd152, 32'sd1501, 32'sd1337, 32'sd1170, 32'sd1034,
32'sd363, 32'sd1808, 32'sd1911, 32'sd1282, 32'sd1814, 32'sd550,
32'sd1643, 32'sd105, 32'sd829, 32'sd814, 32'sd1102, 32'sd1581,
32'sd1296, 32'sd740, 32'sd1581, 32'sd130, 32'sd1433, 32'sd544,
32'sd1777, 32'sd1577, 32'sd1796, 32'sd1178, 32'sd1632, 32'sd1377,
32'sd861, 32'sd1834, 32'sd1859, 32'sd1226, 32'sd1496, 32'sd355,
32'sd1119, 32'sd1979, 32'sd534, 32'sd822, 32'sd388, 32'sd979,
32'sd545, 32'sd1693, 32'sd342, 32'sd627, 32'sd852, 32'sd1030,
32'sd1399, 32'sd1368, 32'sd1775, 32'sd559, 32'sd772, 32'sd1329,
32'sd1900, 32'sd605, 32'sd1801, 32'sd650, 32'sd1924, 32'sd907,
32'sd767, 32'sd1594, 32'sd1247, 32'sd1244, 32'sd782, 32'sd1290,
32'sd1047, 32'sd792, 32'sd1257, 32'sd1273, 32'sd553, 32'sd1711,
32'sd131, 32'sd1907, 32'sd1071, 32'sd407, 32'sd414, 32'sd1392,
32'sd397, 32'sd1274, 32'sd1767, 32'sd687, 32'sd1234, 32'sd1954,
32'sd1594, 32'sd1625, 32'sd1374, 32'sd1211, 32'sd734, 32'sd1133,
32'sd420, 32'sd1685, 32'sd1019, 32'sd237, 32'sd1720, 32'sd1066,
32'sd1626, 32'sd680, 32'sd1542, 32'sd865, 32'sd1342, 32'sd656,
32'sd925, 32'sd856, 32'sd1252, 32'sd1265, 32'sd1730, 32'sd1888,
32'sd1358, 32'sd1089, 32'sd147, 32'sd782, 32'sd1825, 32'sd1773,
32'sd890, 32'sd1397, 32'sd1623, 32'sd1591, 32'sd1027, 32'sd383,
32'sd1918, 32'sd160, 32'sd407, 32'sd224, 32'sd954, 32'sd1440,
32'sd1580, 32'sd213, 32'sd862, 32'sd1054, 32'sd422, 32'sd1459,
32'sd690, 32'sd962, 32'sd1047, 32'sd1524, 32'sd144, 32'sd915,
32'sd1704, 32'sd768, 32'sd159, 32'sd820, 32'sd1294, 32'sd1658,
32'sd525, 32'sd1761, 32'sd1376, 32'sd225, 32'sd748, 32'sd617,
32'sd1127, 32'sd1116, 32'sd1120, 32'sd1259, 32'sd842, 32'sd1829,
32'sd909, 32'sd1634, 32'sd1413, 32'sd1782, 32'sd340, 32'sd1656,
32'sd159, 32'sd874, 32'sd1024, 32'sd1822, 32'sd445, 32'sd952,
32'sd177, 32'sd1593, 32'sd129, 32'sd1027, 32'sd664, 32'sd1208,
32'sd508, 32'sd304, 32'sd1934, 32'sd353, 32'sd670, 32'sd1259,
32'sd219, 32'sd802, 32'sd349, 32'sd1607, 32'sd1125, 32'sd819,
32'sd1538, 32'sd1933, 32'sd455, 32'sd887, 32'sd279, 32'sd1387,
32'sd986, 32'sd271, 32'sd1624, 32'sd1664, 32'sd1362, 32'sd526,
32'sd1655, 32'sd1621, 32'sd907, 32'sd1468, 32'sd1447, 32'sd188,
32'sd281, 32'sd566, 32'sd1404, 32'sd1433, 32'sd1624, 32'sd1580,
32'sd877, 32'sd488, 32'sd355, 32'sd485, 32'sd493, 32'sd1945,
32'sd1000, 32'sd961, 32'sd711, 32'sd697, 32'sd527, 32'sd162,
32'sd1265, 32'sd123, 32'sd1899, 32'sd1287, 32'sd1144, 32'sd1885,
32'sd1453, 32'sd1191, 32'sd243, 32'sd1751, 32'sd840, 32'sd214,
32'sd1784, 32'sd252, 32'sd214, 32'sd642, 32'sd1539, 32'sd605,
32'sd1692, 32'sd466, 32'sd1147, 32'sd737, 32'sd1704, 32'sd1582,
32'sd1056, 32'sd337, 32'sd1683, 32'sd1037, 32'sd519, 32'sd1751,
32'sd263, 32'sd679, 32'sd977, 32'sd1749, 32'sd130, 32'sd1779,
32'sd299, 32'sd624, 32'sd1175, 32'sd1998, 32'sd1154, 32'sd1022,
32'sd274, 32'sd1067, 32'sd1164, 32'sd635, 32'sd252, 32'sd1462,
32'sd183, 32'sd1535, 32'sd375, 32'sd410, 32'sd952, 32'sd1633,
32'sd100, 32'sd930, 32'sd1781, 32'sd598, 32'sd1999, 32'sd266,
32'sd1872, 32'sd1177, 32'sd1627, 32'sd1214, 32'sd1338, 32'sd328,
32'sd1020, 32'sd1164, 32'sd917, 32'sd1665, 32'sd750, 32'sd1222,
32'sd716, 32'sd663, 32'sd1575, 32'sd1886, 32'sd1971, 32'sd1162,
32'sd1008, 32'sd1914, 32'sd859, 32'sd960, 32'sd1454, 32'sd1029,
32'sd977, 32'sd492, 32'sd1506, 32'sd131, 32'sd171, 32'sd1306,
32'sd597, 32'sd688, 32'sd832, 32'sd1224, 32'sd1057, 32'sd1206,
32'sd634, 32'sd1191, 32'sd1019, 32'sd1867, 32'sd647, 32'sd653,
32'sd1668, 32'sd410, 32'sd1228, 32'sd973, 32'sd282, 32'sd100,
32'sd461, 32'sd1507, 32'sd1600, 32'sd1423, 32'sd1618, 32'sd1893,
32'sd954, 32'sd1288, 32'sd125, 32'sd1709, 32'sd363, 32'sd680,
32'sd168, 32'sd347, 32'sd518, 32'sd240, 32'sd938, 32'sd1893,
32'sd1099, 32'sd1983, 32'sd1825, 32'sd1381, 32'sd579, 32'sd586,
32'sd612, 32'sd1189, 32'sd1881, 32'sd466, 32'sd1678, 32'sd1727,
32'sd1539, 32'sd1565, 32'sd524, 32'sd1491, 32'sd706, 32'sd727,
32'sd1423, 32'sd1310, 32'sd1591, 32'sd1296, 32'sd675, 32'sd680,
32'sd800, 32'sd123, 32'sd1259, 32'sd1156, 32'sd436, 32'sd1890,
32'sd1184, 32'sd1601, 32'sd931, 32'sd1295, 32'sd1947, 32'sd1353,
32'sd962, 32'sd887, 32'sd388, 32'sd1611, 32'sd150, 32'sd1732,
32'sd532, 32'sd1427, 32'sd1307, 32'sd1398, 32'sd1176, 32'sd1959,
32'sd589, 32'sd625, 32'sd360, 32'sd1506, 32'sd1076, 32'sd381,
32'sd1061, 32'sd751, 32'sd608, 32'sd1427, 32'sd1293, 32'sd1334,
32'sd230, 32'sd1601, 32'sd1264, 32'sd1953, 32'sd1430, 32'sd1614,
32'sd1778, 32'sd691, 32'sd1347, 32'sd746, 32'sd1237, 32'sd1690,
32'sd1397, 32'sd1011, 32'sd290, 32'sd539, 32'sd335, 32'sd1897,
32'sd201, 32'sd440, 32'sd1897, 32'sd1356, 32'sd855, 32'sd297,
32'sd1917, 32'sd1788, 32'sd1468, 32'sd1903, 32'sd1483, 32'sd1898,
32'sd852, 32'sd1901, 32'sd1544, 32'sd1051, 32'sd1817, 32'sd904,
32'sd648, 32'sd634, 32'sd1267, 32'sd240, 32'sd475, 32'sd739,
32'sd1406, 32'sd1136, 32'sd341, 32'sd1748, 32'sd1602, 32'sd760,
32'sd679, 32'sd1370, 32'sd261, 32'sd1509, 32'sd1782, 32'sd910,
32'sd1345, 32'sd1472, 32'sd1531, 32'sd396, 32'sd936, 32'sd523,
32'sd774, 32'sd703, 32'sd1410, 32'sd862, 32'sd395, 32'sd739,
32'sd1672, 32'sd1608, 32'sd837, 32'sd822, 32'sd370, 32'sd401,
32'sd1802, 32'sd1531, 32'sd1581, 32'sd1018, 32'sd592, 32'sd374,
32'sd125, 32'sd454, 32'sd917, 32'sd1468, 32'sd1321, 32'sd1864,
32'sd416, 32'sd1451, 32'sd1039, 32'sd1859, 32'sd1212, 32'sd206,
32'sd564, 32'sd249, 32'sd922, 32'sd116, 32'sd882, 32'sd323,
32'sd458, 32'sd1554, 32'sd1848, 32'sd1204, 32'sd612, 32'sd1296,
32'sd309, 32'sd998, 32'sd1998, 32'sd1484, 32'sd1731, 32'sd782,
32'sd1320, 32'sd211, 32'sd1113, 32'sd500, 32'sd1216, 32'sd1780,
32'sd1429, 32'sd1119, 32'sd797, 32'sd1607, 32'sd1110, 32'sd1284,
32'sd1989, 32'sd1117, 32'sd480, 32'sd1653, 32'sd107, 32'sd377,
32'sd1918, 32'sd328, 32'sd606, 32'sd1586, 32'sd1411, 32'sd1932,
32'sd332, 32'sd639, 32'sd1062, 32'sd136, 32'sd301, 32'sd721,
32'sd1816, 32'sd863, 32'sd819, 32'sd741, 32'sd246, 32'sd1672,
32'sd1160, 32'sd1428, 32'sd1274, 32'sd107, 32'sd1815, 32'sd1647,
32'sd1175, 32'sd583, 32'sd1806, 32'sd739, 32'sd660, 32'sd1610,
32'sd967, 32'sd123, 32'sd1814, 32'sd102, 32'sd1693, 32'sd193,
32'sd525, 32'sd221, 32'sd1684, 32'sd236, 32'sd549, 32'sd280,
32'sd126, 32'sd889, 32'sd180, 32'sd891, 32'sd688, 32'sd358,
32'sd359, 32'sd523, 32'sd1876, 32'sd166, 32'sd1638, 32'sd1285,
32'sd292, 32'sd1574, 32'sd808, 32'sd434, 32'sd1617, 32'sd345,
32'sd1871, 32'sd622, 32'sd1317, 32'sd983, 32'sd1108, 32'sd1821,
32'sd647, 32'sd1261, 32'sd1157, 32'sd214, 32'sd1310, 32'sd1918,
32'sd1312, 32'sd1040, 32'sd1552, 32'sd1345, 32'sd406, 32'sd1551,
32'sd1748, 32'sd599, 32'sd1163, 32'sd872, 32'sd682, 32'sd1804,
32'sd784, 32'sd1934, 32'sd479, 32'sd402, 32'sd1447, 32'sd1355,
32'sd841, 32'sd1050, 32'sd1177, 32'sd1071, 32'sd1895, 32'sd921,
32'sd133, 32'sd110, 32'sd780, 32'sd1690, 32'sd753, 32'sd145,
32'sd1191, 32'sd222, 32'sd1680, 32'sd1858, 32'sd1788, 32'sd627,
32'sd1196, 32'sd1151, 32'sd267, 32'sd1907, 32'sd152, 32'sd1499,
32'sd1736, 32'sd1041, 32'sd1509, 32'sd1136, 32'sd1256, 32'sd863,
32'sd1322, 32'sd1998, 32'sd1224, 32'sd917, 32'sd1391, 32'sd1736,
32'sd1390, 32'sd561, 32'sd1703, 32'sd1551, 32'sd1042, 32'sd781,
32'sd466, 32'sd1879, 32'sd815, 32'sd1103, 32'sd199, 32'sd216,
32'sd713, 32'sd1884, 32'sd1851, 32'sd215, 32'sd722, 32'sd1722,
32'sd1436, 32'sd1285, 32'sd144, 32'sd1445, 32'sd534, 32'sd1341,
32'sd636, 32'sd1063, 32'sd766, 32'sd207, 32'sd1546, 32'sd1261,
32'sd1185, 32'sd901, 32'sd115, 32'sd892, 32'sd1530, 32'sd1858,
32'sd653, 32'sd510, 32'sd1322, 32'sd900, 32'sd855, 32'sd1845,
32'sd185, 32'sd1095, 32'sd542, 32'sd1674, 32'sd1812, 32'sd164,
32'sd457, 32'sd134, 32'sd509, 32'sd642, 32'sd1977, 32'sd1452,
32'sd742, 32'sd875, 32'sd1075, 32'sd434, 32'sd1649, 32'sd1340,
32'sd1361, 32'sd1318, 32'sd1489, 32'sd468, 32'sd1695, 32'sd1778,
32'sd672, 32'sd1369, 32'sd1960, 32'sd1401, 32'sd165, 32'sd1600,
32'sd1522, 32'sd221, 32'sd1007, 32'sd1984, 32'sd1585, 32'sd963,
32'sd986, 32'sd1566, 32'sd1963, 32'sd1190, 32'sd1527, 32'sd1982,
32'sd934, 32'sd1999, 32'sd1758, 32'sd476, 32'sd1488, 32'sd1112,
32'sd1936, 32'sd529, 32'sd1716, 32'sd1434, 32'sd285, 32'sd1914,
32'sd469, 32'sd725, 32'sd806, 32'sd714, 32'sd451, 32'sd894,
32'sd1052, 32'sd812, 32'sd597, 32'sd729, 32'sd440, 32'sd1546,
32'sd131, 32'sd420, 32'sd1229, 32'sd1377, 32'sd851, 32'sd1564,
32'sd560, 32'sd257, 32'sd968, 32'sd780, 32'sd1114, 32'sd509,
32'sd681, 32'sd564, 32'sd207, 32'sd1619, 32'sd1196, 32'sd542,
32'sd871, 32'sd1358, 32'sd504, 32'sd799, 32'sd563, 32'sd1460,
32'sd1593, 32'sd206, 32'sd1061, 32'sd898, 32'sd868, 32'sd1039,
32'sd1850, 32'sd1387, 32'sd1136, 32'sd150, 32'sd1954, 32'sd1961,
32'sd294, 32'sd1142, 32'sd1586, 32'sd724, 32'sd785, 32'sd1247,
32'sd1349, 32'sd1281, 32'sd799, 32'sd1348, 32'sd1793, 32'sd1205,
32'sd613, 32'sd795, 32'sd1172, 32'sd1317, 32'sd1032, 32'sd1595,
32'sd1173, 32'sd711, 32'sd1792, 32'sd310, 32'sd269, 32'sd1461,
32'sd1635, 32'sd1551, 32'sd792, 32'sd1756, 32'sd1001, 32'sd1278,
32'sd597, 32'sd1084, 32'sd1890, 32'sd1292, 32'sd198, 32'sd597,
32'sd463, 32'sd1551, 32'sd542, 32'sd1151, 32'sd329, 32'sd434,
32'sd1782, 32'sd1344, 32'sd918, 32'sd801, 32'sd1688, 32'sd1911,
32'sd1977, 32'sd404, 32'sd1352, 32'sd489, 32'sd944, 32'sd972,
32'sd1055, 32'sd899, 32'sd573, 32'sd1657, 32'sd939, 32'sd1782,
32'sd898, 32'sd1700, 32'sd1011, 32'sd1456, 32'sd1335, 32'sd1756,
32'sd1605, 32'sd1552, 32'sd1587, 32'sd581, 32'sd662, 32'sd292,
32'sd1507, 32'sd328, 32'sd1669, 32'sd1684, 32'sd1881, 32'sd385,
32'sd608, 32'sd626, 32'sd802, 32'sd851, 32'sd1694, 32'sd767,
32'sd821, 32'sd1141, 32'sd1098, 32'sd1799, 32'sd852, 32'sd722,
32'sd367, 32'sd494, 32'sd601, 32'sd1644, 32'sd1714, 32'sd1540,
32'sd1616, 32'sd992, 32'sd1913, 32'sd336, 32'sd870, 32'sd1731,
32'sd417, 32'sd331, 32'sd833, 32'sd908, 32'sd1076, 32'sd371,
32'sd829, 32'sd1605, 32'sd331, 32'sd1592, 32'sd1913, 32'sd1550,
32'sd956, 32'sd1507, 32'sd568, 32'sd1260, 32'sd1132, 32'sd1725,
32'sd1319, 32'sd1465, 32'sd156, 32'sd1241, 32'sd1827, 32'sd1071,
32'sd1258, 32'sd1424, 32'sd1106, 32'sd416, 32'sd233, 32'sd1696,
32'sd1897, 32'sd2000, 32'sd1434, 32'sd1975, 32'sd1705, 32'sd1220,
32'sd1535, 32'sd780, 32'sd126, 32'sd1977, 32'sd390, 32'sd1518,
32'sd1183, 32'sd337, 32'sd681, 32'sd1838, 32'sd129, 32'sd701,
32'sd1489, 32'sd770, 32'sd1165, 32'sd311, 32'sd444, 32'sd602,
32'sd1378, 32'sd1639, 32'sd1284, 32'sd1729, 32'sd1459, 32'sd377,
32'sd1044, 32'sd1971, 32'sd1757, 32'sd1557, 32'sd1072, 32'sd1596,
32'sd1436, 32'sd1853, 32'sd770, 32'sd1093, 32'sd1405, 32'sd1244,
32'sd1025, 32'sd1329, 32'sd312, 32'sd1562, 32'sd602, 32'sd218,
32'sd1642, 32'sd415, 32'sd1765, 32'sd368, 32'sd849, 32'sd533,
32'sd1639, 32'sd1783, 32'sd1854, 32'sd1109, 32'sd1784, 32'sd1656,
32'sd1971, 32'sd1264, 32'sd1700, 32'sd1734, 32'sd813, 32'sd1692,
32'sd547, 32'sd1276, 32'sd518, 32'sd1376, 32'sd458, 32'sd393,
32'sd602, 32'sd824, 32'sd1869, 32'sd1771, 32'sd833, 32'sd579,
32'sd884, 32'sd1223, 32'sd730, 32'sd1327, 32'sd681, 32'sd1158,
32'sd737, 32'sd856, 32'sd888, 32'sd1342, 32'sd801, 32'sd375,
32'sd566, 32'sd1571, 32'sd540, 32'sd1244, 32'sd1384, 32'sd1718,
32'sd1962, 32'sd288, 32'sd348, 32'sd1521, 32'sd436, 32'sd1795,
32'sd878, 32'sd1519, 32'sd1566, 32'sd1480, 32'sd124, 32'sd1474,
32'sd859, 32'sd298, 32'sd1858, 32'sd872, 32'sd1882, 32'sd991,
32'sd1073, 32'sd783, 32'sd1868, 32'sd105, 32'sd1432, 32'sd665,
32'sd914, 32'sd1153, 32'sd966, 32'sd426, 32'sd291, 32'sd1125,
32'sd1037, 32'sd1825, 32'sd690, 32'sd930, 32'sd1785, 32'sd1049,
32'sd759, 32'sd860, 32'sd1316, 32'sd1250, 32'sd450, 32'sd689,
32'sd588, 32'sd893, 32'sd1943, 32'sd627, 32'sd536, 32'sd1705,
32'sd194, 32'sd977, 32'sd852, 32'sd1612, 32'sd1737, 32'sd1781,
32'sd1754, 32'sd221, 32'sd1210, 32'sd619, 32'sd860, 32'sd1133,
32'sd1261, 32'sd1215, 32'sd552, 32'sd1846, 32'sd322, 32'sd905,
32'sd1437, 32'sd1597, 32'sd735, 32'sd907, 32'sd478, 32'sd1550,
32'sd1000, 32'sd694, 32'sd120, 32'sd1686, 32'sd448, 32'sd984,
32'sd546, 32'sd1179, 32'sd516, 32'sd262, 32'sd1037, 32'sd1423,
32'sd1010, 32'sd1560, 32'sd962, 32'sd1610, 32'sd1848, 32'sd1607,
32'sd1522, 32'sd1074, 32'sd510, 32'sd1377, 32'sd1448, 32'sd557,
32'sd664, 32'sd1237, 32'sd1669, 32'sd1599, 32'sd762, 32'sd334,
32'sd1730, 32'sd1305, 32'sd1726, 32'sd1146, 32'sd1490, 32'sd1175,
32'sd1654, 32'sd388, 32'sd1317, 32'sd1447, 32'sd936, 32'sd421,
32'sd921, 32'sd966, 32'sd881, 32'sd827, 32'sd1902, 32'sd1899,
32'sd1647, 32'sd1891, 32'sd1221, 32'sd1050, 32'sd267, 32'sd1840,
32'sd606, 32'sd941, 32'sd1308, 32'sd1024, 32'sd1735, 32'sd594,
32'sd1362, 32'sd1090, 32'sd113, 32'sd1875, 32'sd1711, 32'sd999,
32'sd1124, 32'sd1759, 32'sd1086, 32'sd536, 32'sd1538, 32'sd988,
32'sd899, 32'sd1703, 32'sd675, 32'sd1569, 32'sd212, 32'sd583,
32'sd111, 32'sd475, 32'sd1346, 32'sd260, 32'sd891, 32'sd819,
32'sd719, 32'sd1449, 32'sd454, 32'sd567, 32'sd717, 32'sd604,
32'sd669, 32'sd827, 32'sd763, 32'sd386, 32'sd1891, 32'sd196,
32'sd650, 32'sd1819, 32'sd1702, 32'sd1584, 32'sd1707, 32'sd534,
32'sd394, 32'sd346, 32'sd820, 32'sd1239, 32'sd491, 32'sd1319,
32'sd377, 32'sd145, 32'sd1286, 32'sd636, 32'sd1522, 32'sd1384,
32'sd1081, 32'sd1196, 32'sd540, 32'sd425, 32'sd1343, 32'sd126,
32'sd538, 32'sd105, 32'sd1357, 32'sd552, 32'sd1743, 32'sd1706,
32'sd497, 32'sd1725, 32'sd1939, 32'sd1623, 32'sd1381, 32'sd1885,
32'sd1686, 32'sd537, 32'sd1183, 32'sd1099, 32'sd283, 32'sd1094,
32'sd278, 32'sd1324, 32'sd257, 32'sd705, 32'sd416, 32'sd1007,
32'sd790, 32'sd1663, 32'sd744, 32'sd702, 32'sd1472, 32'sd1331,
32'sd1580, 32'sd1083, 32'sd187, 32'sd1710, 32'sd614, 32'sd838,
32'sd357, 32'sd1226, 32'sd713, 32'sd1575, 32'sd992, 32'sd898,
32'sd1413, 32'sd1791, 32'sd491, 32'sd462, 32'sd866, 32'sd399,
32'sd1470, 32'sd128, 32'sd1267, 32'sd1386, 32'sd1591, 32'sd854,
32'sd1998, 32'sd1947, 32'sd936, 32'sd789, 32'sd1998, 32'sd1969,
32'sd1799, 32'sd871, 32'sd1239, 32'sd777, 32'sd1996, 32'sd1299,
32'sd1771, 32'sd1529, 32'sd971, 32'sd997, 32'sd247, 32'sd1061,
32'sd602, 32'sd1242, 32'sd1109, 32'sd1727, 32'sd350, 32'sd1558,
32'sd1903, 32'sd461, 32'sd1958, 32'sd1447, 32'sd482, 32'sd1490,
32'sd500, 32'sd1126, 32'sd951, 32'sd844, 32'sd1266, 32'sd698,
32'sd300, 32'sd111, 32'sd1569, 32'sd1485, 32'sd1378, 32'sd553,
32'sd1123, 32'sd711, 32'sd862, 32'sd1031, 32'sd458, 32'sd1024,
32'sd1644, 32'sd262, 32'sd583, 32'sd1220, 32'sd1027, 32'sd1828,
32'sd1882, 32'sd1932, 32'sd918, 32'sd1691, 32'sd1856, 32'sd626,
32'sd948, 32'sd700, 32'sd1719, 32'sd335, 32'sd613, 32'sd892,
32'sd1311, 32'sd930, 32'sd339, 32'sd691, 32'sd1963, 32'sd966,
32'sd1527, 32'sd1074, 32'sd236, 32'sd1262, 32'sd1008, 32'sd1824,
32'sd1950, 32'sd1816, 32'sd309, 32'sd1933, 32'sd592, 32'sd772,
32'sd1699, 32'sd196, 32'sd1244, 32'sd1103, 32'sd964, 32'sd221,
32'sd349, 32'sd130, 32'sd1782, 32'sd148, 32'sd658, 32'sd1225,
32'sd466, 32'sd1731, 32'sd1124, 32'sd325, 32'sd1409, 32'sd992,
32'sd1717, 32'sd1793, 32'sd890, 32'sd608, 32'sd864, 32'sd1078,
32'sd1731, 32'sd1935, 32'sd423, 32'sd380, 32'sd892, 32'sd711,
32'sd1013, 32'sd1999, 32'sd1051, 32'sd1513, 32'sd300, 32'sd1121,
32'sd262, 32'sd1818, 32'sd1138, 32'sd908, 32'sd1448, 32'sd374,
32'sd1712, 32'sd1649, 32'sd492, 32'sd1023, 32'sd935, 32'sd1483,
32'sd1483, 32'sd402, 32'sd1602, 32'sd1313, 32'sd1600, 32'sd496,
32'sd1877, 32'sd575, 32'sd1684, 32'sd1487, 32'sd438, 32'sd1913,
32'sd1618, 32'sd1486, 32'sd1842, 32'sd1954, 32'sd1247, 32'sd1811,
32'sd1309, 32'sd1231, 32'sd1341, 32'sd1206, 32'sd113, 32'sd973,
32'sd490, 32'sd365, 32'sd778, 32'sd1996, 32'sd662, 32'sd1323,
32'sd1604, 32'sd1236, 32'sd267, 32'sd1563, 32'sd1114, 32'sd419,
32'sd1674, 32'sd1582, 32'sd186, 32'sd603, 32'sd520, 32'sd1612,
32'sd1555, 32'sd1810, 32'sd1664, 32'sd809, 32'sd281, 32'sd1118,
32'sd1644, 32'sd1281, 32'sd747, 32'sd679, 32'sd780, 32'sd234,
32'sd1168, 32'sd801, 32'sd1901, 32'sd373, 32'sd761, 32'sd1623,
32'sd1398, 32'sd324, 32'sd1242, 32'sd486, 32'sd1483, 32'sd1840,
32'sd336, 32'sd577, 32'sd990, 32'sd1279, 32'sd1211, 32'sd1265,
32'sd523, 32'sd664, 32'sd1602, 32'sd1105, 32'sd1736, 32'sd1669,
32'sd839, 32'sd1594, 32'sd165, 32'sd1878, 32'sd1822, 32'sd1816,
32'sd930, 32'sd1636, 32'sd1234, 32'sd1820, 32'sd1528, 32'sd1642,
32'sd360, 32'sd1204, 32'sd1238, 32'sd1725, 32'sd905, 32'sd525,
32'sd1930, 32'sd672, 32'sd1398, 32'sd849, 32'sd1569, 32'sd1395,
32'sd1639, 32'sd1591, 32'sd791, 32'sd963, 32'sd1270, 32'sd1084,
32'sd1771, 32'sd704, 32'sd1256, 32'sd590, 32'sd1579, 32'sd1724,
32'sd1510, 32'sd1859, 32'sd1155, 32'sd1721, 32'sd804, 32'sd263,
32'sd1249, 32'sd1977, 32'sd1086, 32'sd885, 32'sd1512, 32'sd1183,
32'sd630, 32'sd1782, 32'sd297, 32'sd1411, 32'sd907, 32'sd1416,
32'sd942, 32'sd614, 32'sd1303, 32'sd681, 32'sd1550, 32'sd1329,
32'sd243, 32'sd1742, 32'sd1271, 32'sd809, 32'sd877, 32'sd476,
32'sd617, 32'sd552, 32'sd716, 32'sd997, 32'sd1477, 32'sd199,
32'sd1088, 32'sd1988, 32'sd781, 32'sd1823, 32'sd973, 32'sd211,
32'sd1180, 32'sd1213, 32'sd1513, 32'sd1976, 32'sd1150, 32'sd896,
32'sd119, 32'sd322, 32'sd868, 32'sd624, 32'sd216, 32'sd543,
32'sd785, 32'sd421, 32'sd1400, 32'sd542, 32'sd771, 32'sd325,
32'sd1750, 32'sd1073, 32'sd548, 32'sd1338, 32'sd472, 32'sd746,
32'sd392, 32'sd494, 32'sd1562, 32'sd1014, 32'sd387, 32'sd544,
32'sd726, 32'sd417, 32'sd1920, 32'sd1489, 32'sd652, 32'sd956,
32'sd445, 32'sd912, 32'sd919, 32'sd133, 32'sd705, 32'sd1502,
32'sd1398, 32'sd1967, 32'sd1090, 32'sd678, 32'sd399, 32'sd1390,
32'sd900, 32'sd747, 32'sd1521, 32'sd1706, 32'sd879, 32'sd1706,
32'sd653, 32'sd1767, 32'sd1901, 32'sd1975, 32'sd736, 32'sd1249,
32'sd1328, 32'sd1704, 32'sd241, 32'sd1372, 32'sd1057, 32'sd1677,
32'sd1615, 32'sd145, 32'sd1149, 32'sd365, 32'sd1611, 32'sd399,
32'sd775, 32'sd658, 32'sd1462, 32'sd1735, 32'sd1724, 32'sd943,
32'sd564, 32'sd325, 32'sd293, 32'sd1646, 32'sd1978, 32'sd257,
32'sd785, 32'sd1677, 32'sd495, 32'sd1082, 32'sd890, 32'sd1890,
32'sd1538, 32'sd1652, 32'sd789, 32'sd300, 32'sd506, 32'sd595,
32'sd431, 32'sd1580, 32'sd1912, 32'sd1882, 32'sd1769, 32'sd171,
32'sd698, 32'sd1414, 32'sd633, 32'sd758, 32'sd1661, 32'sd1851,
32'sd631, 32'sd515, 32'sd1303, 32'sd1042, 32'sd1049, 32'sd496,
32'sd518, 32'sd1084, 32'sd343, 32'sd444, 32'sd1043, 32'sd892,
32'sd1503, 32'sd705, 32'sd928, 32'sd948, 32'sd467, 32'sd381,
32'sd1488, 32'sd1147, 32'sd1842, 32'sd1375, 32'sd1423, 32'sd1706,
32'sd1737, 32'sd783, 32'sd244, 32'sd689, 32'sd386, 32'sd1448,
32'sd1407, 32'sd1790, 32'sd1125, 32'sd353, 32'sd1465, 32'sd278,
32'sd847, 32'sd586, 32'sd1094, 32'sd854, 32'sd1097, 32'sd1265,
32'sd1254, 32'sd616, 32'sd957, 32'sd1446, 32'sd157, 32'sd1331,
32'sd1891, 32'sd738, 32'sd1296, 32'sd125, 32'sd1801, 32'sd1055,
32'sd701, 32'sd1345, 32'sd705, 32'sd866, 32'sd583, 32'sd1705,
32'sd446, 32'sd1880, 32'sd494, 32'sd1424, 32'sd450, 32'sd1540,
32'sd1578, 32'sd1887, 32'sd350, 32'sd1972, 32'sd481, 32'sd1895,
32'sd1292, 32'sd448, 32'sd1593, 32'sd1993, 32'sd1454, 32'sd1616,
32'sd945, 32'sd641, 32'sd1305, 32'sd535, 32'sd994, 32'sd1610,
32'sd1734, 32'sd1655, 32'sd1249, 32'sd1014, 32'sd233, 32'sd1279,
32'sd1981, 32'sd332, 32'sd980, 32'sd1418, 32'sd1864, 32'sd1104,
32'sd231, 32'sd960, 32'sd1365, 32'sd507, 32'sd1319, 32'sd807,
32'sd1764, 32'sd573, 32'sd755, 32'sd409, 32'sd238, 32'sd765,
32'sd832, 32'sd1929, 32'sd241, 32'sd1463, 32'sd1055, 32'sd1103,
32'sd1546, 32'sd1267, 32'sd744, 32'sd786, 32'sd351, 32'sd1573,
32'sd1441, 32'sd366, 32'sd1301, 32'sd1295, 32'sd641, 32'sd843,
32'sd426, 32'sd462, 32'sd1074, 32'sd718, 32'sd531, 32'sd1774,
32'sd304, 32'sd505, 32'sd1853, 32'sd415, 32'sd1502, 32'sd334,
32'sd1625, 32'sd586, 32'sd1611, 32'sd970, 32'sd1649, 32'sd1967,
32'sd1907, 32'sd1449, 32'sd888, 32'sd146, 32'sd1033, 32'sd208,
32'sd467, 32'sd1267, 32'sd265, 32'sd1048, 32'sd893, 32'sd1419,
32'sd1412, 32'sd276, 32'sd256, 32'sd646, 32'sd1482, 32'sd1980,
32'sd923, 32'sd886, 32'sd1195, 32'sd679, 32'sd482, 32'sd1054,
32'sd1689, 32'sd828, 32'sd1622, 32'sd444, 32'sd358, 32'sd517,
32'sd1754, 32'sd1593, 32'sd167, 32'sd216, 32'sd1503, 32'sd101,
32'sd412, 32'sd654, 32'sd681, 32'sd666, 32'sd489, 32'sd681,
32'sd711, 32'sd910, 32'sd472, 32'sd1714, 32'sd1813, 32'sd616,
32'sd647, 32'sd1644, 32'sd1047, 32'sd578, 32'sd280, 32'sd706,
32'sd1078, 32'sd476, 32'sd1807, 32'sd1641, 32'sd1991, 32'sd607,
32'sd1086, 32'sd1689, 32'sd1292, 32'sd332, 32'sd665, 32'sd1781,
32'sd1696, 32'sd1121, 32'sd1875, 32'sd1303, 32'sd609, 32'sd1038,
32'sd1902, 32'sd146, 32'sd541, 32'sd1099, 32'sd1870, 32'sd1607,
32'sd1084, 32'sd222, 32'sd428, 32'sd881, 32'sd245, 32'sd506,
32'sd1300, 32'sd592, 32'sd1928, 32'sd657, 32'sd1032, 32'sd766,
32'sd1564, 32'sd956, 32'sd673, 32'sd1126, 32'sd1701, 32'sd1136,
32'sd933, 32'sd1811, 32'sd1787, 32'sd1400, 32'sd135, 32'sd973,
32'sd696, 32'sd1874, 32'sd1024, 32'sd1914, 32'sd552, 32'sd1167,
32'sd160, 32'sd1325, 32'sd1921, 32'sd1956, 32'sd264, 32'sd887,
32'sd627, 32'sd140, 32'sd1528, 32'sd590, 32'sd1305, 32'sd557,
32'sd1051, 32'sd1816, 32'sd1802, 32'sd108, 32'sd1584, 32'sd1159,
32'sd261, 32'sd721, 32'sd888, 32'sd139, 32'sd1165, 32'sd789,
32'sd348, 32'sd873, 32'sd1388, 32'sd361, 32'sd1900, 32'sd1639,
32'sd1036, 32'sd182, 32'sd1150, 32'sd1687, 32'sd335, 32'sd359,
32'sd902, 32'sd1442, 32'sd1594, 32'sd1239, 32'sd693, 32'sd852,
32'sd1238, 32'sd1535, 32'sd726, 32'sd532, 32'sd1585, 32'sd635,
32'sd1054, 32'sd1366, 32'sd1576, 32'sd996, 32'sd298, 32'sd922,
32'sd698, 32'sd1584, 32'sd532, 32'sd1595, 32'sd1972, 32'sd1382,
32'sd1378, 32'sd852, 32'sd1102, 32'sd411, 32'sd606, 32'sd1042,
32'sd874, 32'sd1160, 32'sd1776, 32'sd527, 32'sd542, 32'sd1891,
32'sd1751, 32'sd1082, 32'sd1763, 32'sd1671, 32'sd409, 32'sd594,
32'sd650, 32'sd643, 32'sd383, 32'sd1430, 32'sd862, 32'sd1827,
32'sd1062, 32'sd1118, 32'sd1377, 32'sd1668, 32'sd295, 32'sd1121,
32'sd1909, 32'sd588, 32'sd1384, 32'sd1913, 32'sd1384, 32'sd1577,
32'sd1638, 32'sd1851, 32'sd952, 32'sd243, 32'sd1953, 32'sd668,
32'sd1648, 32'sd550, 32'sd1668, 32'sd1590, 32'sd943, 32'sd1845,
32'sd1896, 32'sd407, 32'sd794, 32'sd1605, 32'sd1595, 32'sd1868,
32'sd987, 32'sd715, 32'sd188, 32'sd1416, 32'sd1418, 32'sd1845,
32'sd1991, 32'sd817, 32'sd889, 32'sd487, 32'sd1370, 32'sd173,
32'sd1584, 32'sd813, 32'sd970, 32'sd1017, 32'sd633, 32'sd250,
32'sd803, 32'sd356, 32'sd731, 32'sd409, 32'sd1259, 32'sd1584,
32'sd1446, 32'sd596, 32'sd1090, 32'sd281, 32'sd1020, 32'sd441,
32'sd1767, 32'sd1516, 32'sd892, 32'sd1340, 32'sd705, 32'sd983,
32'sd196, 32'sd1610, 32'sd1451, 32'sd1428, 32'sd1442, 32'sd1543,
32'sd989, 32'sd1854, 32'sd1085, 32'sd1426, 32'sd1618, 32'sd1876,
32'sd1408, 32'sd1773, 32'sd685, 32'sd1801, 32'sd238, 32'sd1030,
32'sd990, 32'sd567, 32'sd461, 32'sd1765, 32'sd1845, 32'sd118,
32'sd1998, 32'sd130, 32'sd1805, 32'sd1690, 32'sd1005, 32'sd1699,
32'sd774, 32'sd1018, 32'sd1792, 32'sd821, 32'sd1880, 32'sd514,
32'sd553, 32'sd1603, 32'sd939, 32'sd1056, 32'sd1350, 32'sd700,
32'sd1329, 32'sd235, 32'sd1878, 32'sd169, 32'sd1898, 32'sd1581,
32'sd783, 32'sd1363, 32'sd102, 32'sd114, 32'sd254, 32'sd598,
32'sd933, 32'sd365, 32'sd1887, 32'sd449, 32'sd362, 32'sd201,
32'sd1317, 32'sd1763, 32'sd1341, 32'sd1752, 32'sd416, 32'sd1908,
32'sd917, 32'sd1125, 32'sd730, 32'sd1783, 32'sd542, 32'sd1950,
32'sd1464, 32'sd1518, 32'sd1474, 32'sd1730, 32'sd1696, 32'sd1195,
32'sd319, 32'sd1416, 32'sd289, 32'sd1494, 32'sd1556, 32'sd120,
32'sd579, 32'sd1818, 32'sd546, 32'sd1719, 32'sd1301, 32'sd961,
32'sd630, 32'sd1222, 32'sd1310, 32'sd321, 32'sd1069, 32'sd494,
32'sd1560, 32'sd1885, 32'sd1442, 32'sd737, 32'sd362, 32'sd1360,
32'sd428, 32'sd622, 32'sd167, 32'sd1553, 32'sd1063, 32'sd1206,
32'sd1535, 32'sd597, 32'sd771, 32'sd1151, 32'sd167, 32'sd1116,
32'sd531, 32'sd1373, 32'sd572, 32'sd980, 32'sd1834, 32'sd276,
32'sd1133, 32'sd1860, 32'sd178, 32'sd276, 32'sd1570, 32'sd1358,
32'sd1917, 32'sd184, 32'sd1256, 32'sd620, 32'sd172, 32'sd149,
32'sd984, 32'sd1995, 32'sd917, 32'sd214, 32'sd1269, 32'sd1487,
32'sd1799, 32'sd1664, 32'sd154, 32'sd1843, 32'sd1067, 32'sd1586,
32'sd1934, 32'sd1813, 32'sd1068, 32'sd359, 32'sd340, 32'sd1267,
32'sd1946, 32'sd1210, 32'sd130, 32'sd535, 32'sd1850, 32'sd641,
32'sd613, 32'sd708, 32'sd649, 32'sd681, 32'sd1506, 32'sd807,
32'sd142, 32'sd1134, 32'sd1687, 32'sd1944, 32'sd627, 32'sd1290,
32'sd1255, 32'sd813, 32'sd776, 32'sd1387, 32'sd1966, 32'sd1452,
32'sd470, 32'sd1161, 32'sd1245, 32'sd1539, 32'sd998, 32'sd1193,
32'sd519, 32'sd1630, 32'sd981, 32'sd1865, 32'sd1801, 32'sd773,
32'sd1181, 32'sd759, 32'sd1300, 32'sd1611, 32'sd1491, 32'sd802,
32'sd237, 32'sd1684, 32'sd214, 32'sd1292, 32'sd854, 32'sd701,
32'sd1426, 32'sd1470, 32'sd1998, 32'sd185, 32'sd424, 32'sd168,
32'sd1039, 32'sd347, 32'sd137, 32'sd1762, 32'sd206, 32'sd1523,
32'sd1669, 32'sd1489, 32'sd1759, 32'sd202, 32'sd388, 32'sd499,
32'sd1780, 32'sd324, 32'sd1253, 32'sd516, 32'sd474, 32'sd852,
32'sd126, 32'sd452, 32'sd629, 32'sd780, 32'sd1149, 32'sd256,
32'sd998, 32'sd1531, 32'sd1592, 32'sd1424, 32'sd330, 32'sd1077,
32'sd1602, 32'sd548, 32'sd1377, 32'sd1809, 32'sd892, 32'sd831,
32'sd1337, 32'sd1237, 32'sd1131, 32'sd100, 32'sd299, 32'sd1305,
32'sd226, 32'sd930, 32'sd199, 32'sd186, 32'sd1280, 32'sd331,
32'sd564, 32'sd666, 32'sd1293, 32'sd1276, 32'sd796, 32'sd224,
32'sd151, 32'sd114, 32'sd1307, 32'sd1011, 32'sd1572, 32'sd146,
32'sd1834, 32'sd1031, 32'sd304, 32'sd766, 32'sd1011, 32'sd1102,
32'sd135, 32'sd1385, 32'sd1264, 32'sd1086, 32'sd443, 32'sd1259,
32'sd1679, 32'sd127, 32'sd1199, 32'sd771, 32'sd237, 32'sd1425,
32'sd1546, 32'sd1343, 32'sd220, 32'sd1595, 32'sd542, 32'sd484,
32'sd1216, 32'sd1489, 32'sd142, 32'sd811, 32'sd620, 32'sd203,
32'sd1929, 32'sd1993, 32'sd1523, 32'sd324, 32'sd316, 32'sd657,
32'sd729, 32'sd661, 32'sd312, 32'sd1149, 32'sd701, 32'sd1891,
32'sd1239, 32'sd1466, 32'sd953, 32'sd155, 32'sd1181, 32'sd1413,
32'sd1526, 32'sd1238, 32'sd1836, 32'sd757, 32'sd1641, 32'sd569,
32'sd1332, 32'sd1420, 32'sd1500, 32'sd904, 32'sd297, 32'sd244,
32'sd1274, 32'sd764, 32'sd835, 32'sd683, 32'sd370, 32'sd1832,
32'sd587, 32'sd812, 32'sd163, 32'sd1626, 32'sd1342, 32'sd180,
32'sd1543, 32'sd1765, 32'sd1326, 32'sd648, 32'sd689, 32'sd1593,
32'sd1520, 32'sd450, 32'sd1116, 32'sd891, 32'sd1923, 32'sd844,
32'sd1674, 32'sd1033, 32'sd982, 32'sd389, 32'sd572, 32'sd528,
32'sd1155, 32'sd812, 32'sd1027, 32'sd1078, 32'sd395, 32'sd1866,
32'sd718, 32'sd1197, 32'sd1868, 32'sd935, 32'sd986, 32'sd1100,
32'sd517, 32'sd1957, 32'sd1886, 32'sd1556, 32'sd819, 32'sd1361,
32'sd1386, 32'sd331, 32'sd438, 32'sd214, 32'sd458, 32'sd1725,
32'sd1910, 32'sd812, 32'sd1356, 32'sd416, 32'sd429, 32'sd1507,
32'sd142, 32'sd1145, 32'sd1237, 32'sd349, 32'sd388, 32'sd161,
32'sd1973, 32'sd798, 32'sd760, 32'sd728, 32'sd821, 32'sd460,
32'sd1744, 32'sd1871, 32'sd276, 32'sd860, 32'sd1480, 32'sd1057,
32'sd708, 32'sd1894, 32'sd1351, 32'sd1320, 32'sd1002, 32'sd1967,
32'sd1261, 32'sd426, 32'sd1000, 32'sd1585, 32'sd1592, 32'sd875,
32'sd1002, 32'sd674, 32'sd1467, 32'sd1603, 32'sd640, 32'sd217,
32'sd214, 32'sd1344, 32'sd1223, 32'sd489, 32'sd1110, 32'sd1663,
32'sd839, 32'sd728, 32'sd399, 32'sd1233, 32'sd167, 32'sd1782,
32'sd1824, 32'sd1178, 32'sd1241, 32'sd1335, 32'sd1806, 32'sd1859,
32'sd1364, 32'sd1437, 32'sd825, 32'sd1191, 32'sd428, 32'sd124,
32'sd1746, 32'sd1561, 32'sd175, 32'sd1612, 32'sd1083, 32'sd557,
32'sd1872, 32'sd1980, 32'sd1669, 32'sd285, 32'sd868, 32'sd700,
32'sd654, 32'sd1294, 32'sd781, 32'sd1698, 32'sd1868, 32'sd937,
32'sd381, 32'sd1153, 32'sd1724, 32'sd1326, 32'sd1437, 32'sd234,
32'sd722, 32'sd1665, 32'sd678, 32'sd338, 32'sd372, 32'sd298,
32'sd1756, 32'sd1599, 32'sd253, 32'sd1802, 32'sd1816, 32'sd1744,
32'sd1044, 32'sd686, 32'sd588, 32'sd1818, 32'sd417, 32'sd730,
32'sd1643, 32'sd1043, 32'sd1120, 32'sd471, 32'sd701, 32'sd1292,
32'sd1656, 32'sd535, 32'sd1426, 32'sd1532, 32'sd828, 32'sd1669,
32'sd1024, 32'sd152, 32'sd1880, 32'sd293, 32'sd1423, 32'sd1668,
32'sd1217, 32'sd593, 32'sd1945, 32'sd225, 32'sd282, 32'sd886,
32'sd1189, 32'sd1038, 32'sd871, 32'sd1196, 32'sd890, 32'sd1771,
32'sd1789, 32'sd281, 32'sd1225, 32'sd1317, 32'sd127, 32'sd940,
32'sd1510, 32'sd1083, 32'sd1348, 32'sd688, 32'sd1198, 32'sd1413,
32'sd1435, 32'sd1400, 32'sd159, 32'sd1586, 32'sd299, 32'sd1204,
32'sd1776, 32'sd406, 32'sd545, 32'sd1283, 32'sd1258, 32'sd1163,
32'sd200, 32'sd356, 32'sd1484, 32'sd223, 32'sd1823, 32'sd1371,
32'sd1350, 32'sd1556, 32'sd1889, 32'sd764, 32'sd1508, 32'sd715,
32'sd1269, 32'sd278, 32'sd957, 32'sd171, 32'sd269, 32'sd452,
32'sd1693, 32'sd1834, 32'sd1812, 32'sd681, 32'sd282, 32'sd1903,
32'sd1007, 32'sd468, 32'sd1877, 32'sd377, 32'sd1885, 32'sd306,
32'sd1172, 32'sd1427, 32'sd1998, 32'sd1380, 32'sd488, 32'sd1215,
32'sd1457, 32'sd1516, 32'sd232, 32'sd433, 32'sd1052, 32'sd927,
32'sd597, 32'sd398, 32'sd103, 32'sd1433, 32'sd1472, 32'sd1334,
32'sd361, 32'sd1491, 32'sd1823, 32'sd507, 32'sd1156, 32'sd521,
32'sd489, 32'sd1286, 32'sd1609, 32'sd1899, 32'sd1103, 32'sd486,
32'sd1893, 32'sd768, 32'sd1328, 32'sd1740, 32'sd1322, 32'sd645,
32'sd1105, 32'sd1407, 32'sd1419, 32'sd828, 32'sd414, 32'sd1416,
32'sd1764, 32'sd916, 32'sd347, 32'sd884, 32'sd1026, 32'sd1831,
32'sd1618, 32'sd1446, 32'sd592, 32'sd1376, 32'sd1481, 32'sd1852,
32'sd1413, 32'sd530, 32'sd1731, 32'sd1578, 32'sd457, 32'sd374,
32'sd705, 32'sd1631, 32'sd1403, 32'sd1786, 32'sd197, 32'sd267,
32'sd717, 32'sd1591, 32'sd1526, 32'sd1224, 32'sd593, 32'sd1266,
32'sd614, 32'sd806, 32'sd267, 32'sd1955, 32'sd1798, 32'sd1906,
32'sd1071, 32'sd1527, 32'sd622, 32'sd1302, 32'sd455, 32'sd1638,
32'sd386, 32'sd164, 32'sd1712, 32'sd1827, 32'sd804, 32'sd1107,
32'sd919, 32'sd1216, 32'sd304, 32'sd598, 32'sd1502, 32'sd1491,
32'sd612, 32'sd221, 32'sd625, 32'sd990, 32'sd1972, 32'sd1840,
32'sd1003, 32'sd1404, 32'sd1436, 32'sd1874, 32'sd1153, 32'sd305,
32'sd261, 32'sd209, 32'sd833, 32'sd1204, 32'sd1654, 32'sd214,
32'sd177, 32'sd496, 32'sd550, 32'sd557, 32'sd1642, 32'sd1773,
32'sd1660, 32'sd1617, 32'sd1694, 32'sd1011, 32'sd1826, 32'sd1394,
32'sd1690, 32'sd684, 32'sd255, 32'sd1204, 32'sd1906, 32'sd1005,
32'sd1508, 32'sd1745, 32'sd1029, 32'sd1292, 32'sd178, 32'sd912,
32'sd241, 32'sd129, 32'sd1900, 32'sd1469, 32'sd1137, 32'sd1700,
32'sd244, 32'sd525, 32'sd470, 32'sd424, 32'sd1682, 32'sd1848,
32'sd834, 32'sd1450, 32'sd125, 32'sd1622, 32'sd1045, 32'sd561,
32'sd509, 32'sd414, 32'sd1759, 32'sd1654, 32'sd1965, 32'sd166,
32'sd1272, 32'sd1933, 32'sd1532, 32'sd149, 32'sd911, 32'sd1192,
32'sd1248, 32'sd239, 32'sd1950, 32'sd1497, 32'sd813, 32'sd1021,
32'sd292, 32'sd1377, 32'sd306, 32'sd1458, 32'sd1501, 32'sd1405,
32'sd1675, 32'sd1083, 32'sd747, 32'sd1080, 32'sd1251, 32'sd187,
32'sd554, 32'sd950, 32'sd294, 32'sd1191, 32'sd1598, 32'sd123,
32'sd1717, 32'sd523, 32'sd1859, 32'sd306, 32'sd1276, 32'sd1317,
32'sd636, 32'sd1570, 32'sd1406, 32'sd565, 32'sd1263, 32'sd652,
32'sd733, 32'sd1976, 32'sd303, 32'sd1481, 32'sd1984, 32'sd1815,
32'sd843, 32'sd1931, 32'sd352, 32'sd673, 32'sd589, 32'sd410,
32'sd578, 32'sd1382, 32'sd356, 32'sd287, 32'sd732, 32'sd1618,
32'sd1343, 32'sd1731, 32'sd830, 32'sd1008, 32'sd822, 32'sd741,
32'sd816, 32'sd909, 32'sd1482, 32'sd791, 32'sd1849, 32'sd124,
32'sd328, 32'sd659, 32'sd1859, 32'sd1287, 32'sd1969, 32'sd842,
32'sd793, 32'sd331, 32'sd470, 32'sd445, 32'sd1073, 32'sd1077,
32'sd405, 32'sd661, 32'sd1008, 32'sd1019, 32'sd926, 32'sd258,
32'sd1433, 32'sd1179, 32'sd1900, 32'sd195, 32'sd1280, 32'sd1300,
32'sd908, 32'sd679, 32'sd1258, 32'sd427, 32'sd115, 32'sd1951,
32'sd1245, 32'sd1778, 32'sd1845, 32'sd1277, 32'sd1377, 32'sd1464,
32'sd1032, 32'sd136, 32'sd472, 32'sd591, 32'sd736, 32'sd307,
32'sd1532, 32'sd364, 32'sd1069, 32'sd1379, 32'sd1359, 32'sd488,
32'sd564, 32'sd1886, 32'sd657, 32'sd1202, 32'sd1003, 32'sd1755,
32'sd1262, 32'sd1086, 32'sd339, 32'sd801, 32'sd1639, 32'sd1977,
32'sd1275, 32'sd269, 32'sd434, 32'sd1294, 32'sd1756, 32'sd1030,
32'sd288, 32'sd338, 32'sd1244, 32'sd547, 32'sd457, 32'sd1779,
32'sd1042, 32'sd991, 32'sd1945, 32'sd1834, 32'sd278, 32'sd1001,
32'sd1366, 32'sd431, 32'sd278, 32'sd1054, 32'sd1461, 32'sd1350,
32'sd1308, 32'sd239, 32'sd1472, 32'sd1692, 32'sd465, 32'sd821,
32'sd1596, 32'sd1166, 32'sd175, 32'sd522, 32'sd1124, 32'sd1160,
32'sd525, 32'sd786, 32'sd1570, 32'sd1335, 32'sd1892, 32'sd1270,
32'sd1486, 32'sd1423, 32'sd167, 32'sd1505, 32'sd1966, 32'sd572,
32'sd179, 32'sd946, 32'sd363, 32'sd539, 32'sd930, 32'sd1980,
32'sd280, 32'sd1398, 32'sd1002, 32'sd1401, 32'sd1321, 32'sd619,
32'sd1293, 32'sd369, 32'sd342, 32'sd1967, 32'sd676, 32'sd379,
32'sd325, 32'sd375, 32'sd814, 32'sd1254, 32'sd952, 32'sd335,
32'sd1125, 32'sd1220, 32'sd1949, 32'sd267, 32'sd741, 32'sd1475,
32'sd1296, 32'sd979, 32'sd553, 32'sd886, 32'sd1764, 32'sd1238,
32'sd293, 32'sd1586, 32'sd245, 32'sd770, 32'sd212, 32'sd678,
32'sd309, 32'sd1476, 32'sd1705, 32'sd697, 32'sd1060, 32'sd1766,
32'sd1293, 32'sd1809, 32'sd1905, 32'sd367, 32'sd1677, 32'sd1685,
32'sd610, 32'sd1948, 32'sd1844, 32'sd1948, 32'sd1319, 32'sd1165,
32'sd483, 32'sd211, 32'sd501, 32'sd647, 32'sd1737, 32'sd588,
32'sd844, 32'sd747, 32'sd937, 32'sd973, 32'sd1266, 32'sd1563,
32'sd251, 32'sd580, 32'sd1447, 32'sd505, 32'sd214, 32'sd1680,
32'sd1654, 32'sd1969, 32'sd1486, 32'sd1582, 32'sd1018, 32'sd1601,
32'sd1468, 32'sd573, 32'sd1013, 32'sd681, 32'sd1184, 32'sd1581,
32'sd186, 32'sd1976, 32'sd493, 32'sd540, 32'sd1951, 32'sd736,
32'sd1281, 32'sd1390, 32'sd109, 32'sd1213, 32'sd1731, 32'sd1407,
32'sd177, 32'sd1204, 32'sd341, 32'sd330, 32'sd1166, 32'sd406,
32'sd870, 32'sd1920, 32'sd888, 32'sd1066, 32'sd533, 32'sd1404,
32'sd1224, 32'sd516, 32'sd1223, 32'sd1090, 32'sd821, 32'sd1415,
32'sd374, 32'sd1634, 32'sd1104, 32'sd1730, 32'sd1501, 32'sd270,
32'sd1400, 32'sd655, 32'sd1057, 32'sd1052, 32'sd1162, 32'sd304,
32'sd624, 32'sd189, 32'sd1375, 32'sd1091, 32'sd773, 32'sd1552,
32'sd1407, 32'sd1854, 32'sd505, 32'sd1846, 32'sd1068, 32'sd1688,
32'sd1402, 32'sd394, 32'sd1900, 32'sd881, 32'sd894, 32'sd132,
32'sd1135, 32'sd828, 32'sd960, 32'sd767, 32'sd1781, 32'sd290,
32'sd1939, 32'sd549, 32'sd1240, 32'sd1674, 32'sd969, 32'sd1297,
32'sd702, 32'sd1017, 32'sd815, 32'sd515, 32'sd1506, 32'sd502,
32'sd1235, 32'sd771, 32'sd1815, 32'sd669, 32'sd1736, 32'sd1043,
32'sd1807, 32'sd762, 32'sd618, 32'sd1356, 32'sd1346, 32'sd1077,
32'sd1995, 32'sd170, 32'sd1260, 32'sd386, 32'sd283, 32'sd1652,
32'sd1100, 32'sd1029, 32'sd764, 32'sd1261, 32'sd642, 32'sd706,
32'sd193, 32'sd1668, 32'sd822, 32'sd1736, 32'sd933, 32'sd1505,
32'sd626, 32'sd1413, 32'sd304, 32'sd1690, 32'sd555, 32'sd346,
32'sd589, 32'sd820, 32'sd990, 32'sd1599, 32'sd1980, 32'sd1443,
32'sd1670, 32'sd1589, 32'sd410, 32'sd1776, 32'sd1185, 32'sd268,
32'sd941, 32'sd1380, 32'sd753, 32'sd503, 32'sd1689, 32'sd1227,
32'sd1430, 32'sd669, 32'sd510, 32'sd454, 32'sd472, 32'sd1849,
32'sd1579, 32'sd335, 32'sd1702, 32'sd582, 32'sd566, 32'sd447,
32'sd1918, 32'sd1997, 32'sd1460, 32'sd741, 32'sd416, 32'sd985,
32'sd256, 32'sd789, 32'sd277, 32'sd1295, 32'sd627, 32'sd1568,
32'sd762, 32'sd1603, 32'sd242, 32'sd1952, 32'sd1628, 32'sd1162,
32'sd996, 32'sd1558, 32'sd918, 32'sd1189, 32'sd1291, 32'sd957,
32'sd1589, 32'sd700, 32'sd1861, 32'sd902, 32'sd1486, 32'sd1118,
32'sd1986, 32'sd1539, 32'sd1158, 32'sd834, 32'sd1262, 32'sd1989,
32'sd506, 32'sd997, 32'sd1189, 32'sd221, 32'sd688, 32'sd730,
32'sd271, 32'sd891, 32'sd572, 32'sd547, 32'sd983, 32'sd1276,
32'sd1354, 32'sd221, 32'sd291, 32'sd319, 32'sd756, 32'sd1846,
32'sd1881, 32'sd115, 32'sd1203, 32'sd845, 32'sd1161, 32'sd1176,
32'sd1661, 32'sd1791, 32'sd845, 32'sd277, 32'sd963, 32'sd1563,
32'sd295, 32'sd523, 32'sd285, 32'sd978, 32'sd438, 32'sd1863,
32'sd1019, 32'sd585, 32'sd509, 32'sd556, 32'sd526, 32'sd121,
32'sd1668, 32'sd739, 32'sd678, 32'sd1207, 32'sd637, 32'sd673,
32'sd461, 32'sd251, 32'sd204, 32'sd312, 32'sd1697, 32'sd187,
32'sd125, 32'sd1486, 32'sd1150, 32'sd333, 32'sd1910, 32'sd1013,
32'sd1032, 32'sd1481, 32'sd558, 32'sd287, 32'sd576, 32'sd261,
32'sd568, 32'sd1767, 32'sd1407, 32'sd1667, 32'sd1324, 32'sd243,
32'sd493, 32'sd923, 32'sd854, 32'sd1092, 32'sd608, 32'sd918,
32'sd1071, 32'sd958, 32'sd707, 32'sd1264, 32'sd180, 32'sd1736,
32'sd155, 32'sd941, 32'sd1355, 32'sd878, 32'sd282, 32'sd610,
32'sd1077, 32'sd1711, 32'sd1679, 32'sd1832, 32'sd888, 32'sd457,
32'sd1872, 32'sd1143, 32'sd1355, 32'sd756, 32'sd1657, 32'sd1120,
32'sd612, 32'sd1217, 32'sd135, 32'sd232, 32'sd1951, 32'sd1737,
32'sd264, 32'sd227, 32'sd1173, 32'sd651, 32'sd1156, 32'sd1774,
32'sd1850, 32'sd1408, 32'sd1025, 32'sd325, 32'sd1199, 32'sd574,
32'sd124, 32'sd559, 32'sd1489, 32'sd1476, 32'sd1987, 32'sd706,
32'sd772, 32'sd961, 32'sd554, 32'sd1152, 32'sd1559, 32'sd1192,
32'sd1051, 32'sd1363, 32'sd848, 32'sd845, 32'sd1762, 32'sd1072,
32'sd1386, 32'sd865, 32'sd1411, 32'sd1768, 32'sd1339, 32'sd917,
32'sd415, 32'sd900, 32'sd946, 32'sd1576, 32'sd1369, 32'sd178,
32'sd1904, 32'sd1492, 32'sd1579, 32'sd365, 32'sd1849, 32'sd1445,
32'sd841, 32'sd514, 32'sd816, 32'sd1994, 32'sd1464, 32'sd1094,
32'sd1060, 32'sd1668, 32'sd1677, 32'sd1313, 32'sd1437, 32'sd1216,
32'sd1016, 32'sd562, 32'sd1455, 32'sd1776, 32'sd313, 32'sd1927,
32'sd1264, 32'sd1071, 32'sd1691, 32'sd736, 32'sd297, 32'sd461,
32'sd622, 32'sd1831, 32'sd598, 32'sd142, 32'sd513, 32'sd181,
32'sd1613, 32'sd1284, 32'sd916, 32'sd1476, 32'sd111, 32'sd769,
32'sd1836, 32'sd457, 32'sd409, 32'sd1345, 32'sd1013, 32'sd213,
32'sd295, 32'sd496, 32'sd1352, 32'sd1513, 32'sd1042, 32'sd1196,
32'sd1652, 32'sd1085, 32'sd924, 32'sd109, 32'sd1486, 32'sd670,
32'sd164, 32'sd440, 32'sd1181, 32'sd549, 32'sd151, 32'sd1731,
32'sd604, 32'sd1448, 32'sd1025, 32'sd1361, 32'sd424, 32'sd1046,
32'sd343, 32'sd479, 32'sd882, 32'sd1068, 32'sd191, 32'sd892,
32'sd1317, 32'sd1130, 32'sd121, 32'sd696, 32'sd1159, 32'sd981,
32'sd824, 32'sd597, 32'sd1649, 32'sd1008, 32'sd1908, 32'sd739,
32'sd1813, 32'sd313, 32'sd307, 32'sd1621, 32'sd1015, 32'sd1333,
32'sd1162, 32'sd1020, 32'sd380, 32'sd1012, 32'sd747, 32'sd1770,
32'sd956, 32'sd167, 32'sd1332, 32'sd104, 32'sd121, 32'sd1067,
32'sd482, 32'sd362, 32'sd1883, 32'sd1891, 32'sd143, 32'sd317,
32'sd922, 32'sd963, 32'sd643, 32'sd1053, 32'sd493, 32'sd888,
32'sd1781, 32'sd387, 32'sd1185, 32'sd917, 32'sd614, 32'sd146,
32'sd1114, 32'sd1986, 32'sd1933, 32'sd566, 32'sd1952, 32'sd200,
32'sd1143, 32'sd574, 32'sd799, 32'sd1556, 32'sd833, 32'sd846,
32'sd1472, 32'sd1540, 32'sd649, 32'sd1856, 32'sd179, 32'sd702,
32'sd512, 32'sd283, 32'sd919, 32'sd786, 32'sd1362, 32'sd171,
32'sd652, 32'sd657, 32'sd614, 32'sd314, 32'sd114, 32'sd983,
32'sd1336, 32'sd263, 32'sd458, 32'sd597, 32'sd385, 32'sd410,
32'sd752, 32'sd1818, 32'sd603, 32'sd1861, 32'sd1181, 32'sd1563,
32'sd489, 32'sd1729, 32'sd615, 32'sd1926, 32'sd412, 32'sd1405,
32'sd1332, 32'sd1514, 32'sd856, 32'sd789, 32'sd498, 32'sd426,
32'sd1861, 32'sd744, 32'sd795, 32'sd519, 32'sd816, 32'sd1191,
32'sd184, 32'sd570, 32'sd129, 32'sd773, 32'sd1883, 32'sd1270,
32'sd1303, 32'sd538, 32'sd1405, 32'sd279, 32'sd430, 32'sd503,
32'sd1296, 32'sd1270, 32'sd1069, 32'sd1841, 32'sd1776, 32'sd363,
32'sd803, 32'sd612, 32'sd1074, 32'sd1121, 32'sd860, 32'sd1663,
32'sd945, 32'sd429, 32'sd1942, 32'sd1083, 32'sd1139, 32'sd1751,
32'sd686, 32'sd798, 32'sd1828, 32'sd499, 32'sd1275, 32'sd666,
32'sd248, 32'sd1529, 32'sd286, 32'sd185, 32'sd987, 32'sd1228,
32'sd1247, 32'sd1636, 32'sd1468, 32'sd1129, 32'sd1859, 32'sd614,
32'sd1841, 32'sd225, 32'sd533, 32'sd1955, 32'sd1829, 32'sd1377,
32'sd1321, 32'sd1884, 32'sd411, 32'sd715, 32'sd383, 32'sd628,
32'sd125, 32'sd1246, 32'sd474, 32'sd241, 32'sd850, 32'sd1928,
32'sd189, 32'sd924, 32'sd249, 32'sd1943, 32'sd1167, 32'sd1737,
32'sd500, 32'sd1191, 32'sd665, 32'sd1836, 32'sd967, 32'sd153,
32'sd1796, 32'sd1683, 32'sd455, 32'sd748, 32'sd715, 32'sd552,
32'sd1722, 32'sd179, 32'sd512, 32'sd788, 32'sd1431, 32'sd1044,
32'sd782, 32'sd1061, 32'sd1513, 32'sd999, 32'sd355, 32'sd898,
32'sd1791, 32'sd1689, 32'sd1922, 32'sd1332, 32'sd917, 32'sd1017,
32'sd704, 32'sd101, 32'sd1818, 32'sd1867, 32'sd1212, 32'sd1339,
32'sd1130, 32'sd1927, 32'sd193, 32'sd1879, 32'sd441, 32'sd1497,
32'sd1302, 32'sd575, 32'sd1518, 32'sd1308, 32'sd1034, 32'sd1019,
32'sd1338, 32'sd482, 32'sd632, 32'sd410, 32'sd226, 32'sd595,
32'sd737, 32'sd194, 32'sd770, 32'sd986, 32'sd942, 32'sd1762,
32'sd589, 32'sd1018, 32'sd1984, 32'sd405, 32'sd1421, 32'sd1398,
32'sd922, 32'sd1083, 32'sd1723, 32'sd1382, 32'sd296, 32'sd1508,
32'sd1395, 32'sd141, 32'sd490, 32'sd243, 32'sd300, 32'sd858,
32'sd438, 32'sd913, 32'sd1959, 32'sd735, 32'sd857, 32'sd1152,
32'sd442, 32'sd1524, 32'sd680, 32'sd1925, 32'sd964, 32'sd909,
32'sd1762, 32'sd154, 32'sd1312, 32'sd1097, 32'sd408, 32'sd1130,
32'sd1369, 32'sd108, 32'sd397, 32'sd653, 32'sd1343, 32'sd1016,
32'sd576, 32'sd1199, 32'sd1100, 32'sd760, 32'sd272, 32'sd265,
32'sd1047, 32'sd943, 32'sd231, 32'sd931, 32'sd322, 32'sd521,
32'sd1387, 32'sd1116, 32'sd1597, 32'sd247, 32'sd1750, 32'sd1285,
32'sd188, 32'sd412, 32'sd347, 32'sd106, 32'sd1628, 32'sd1680,
32'sd921, 32'sd727, 32'sd1935, 32'sd1102, 32'sd948, 32'sd386,
32'sd1650, 32'sd967, 32'sd1884, 32'sd727, 32'sd742, 32'sd1124,
32'sd442, 32'sd743, 32'sd1108, 32'sd228, 32'sd853, 32'sd1833,
32'sd1535, 32'sd1485, 32'sd268, 32'sd171, 32'sd1501, 32'sd420,
32'sd100, 32'sd1119, 32'sd1794, 32'sd676, 32'sd617, 32'sd359,
32'sd361, 32'sd458, 32'sd1732, 32'sd141, 32'sd214, 32'sd1094,
32'sd442, 32'sd513, 32'sd1689, 32'sd245, 32'sd313, 32'sd329,
32'sd1277, 32'sd1292, 32'sd122, 32'sd1005, 32'sd1514, 32'sd1132,
32'sd544, 32'sd1298, 32'sd936, 32'sd386, 32'sd1956, 32'sd127,
32'sd608, 32'sd1185, 32'sd870, 32'sd1998, 32'sd1425, 32'sd881,
32'sd1680, 32'sd1351, 32'sd1746, 32'sd463, 32'sd979, 32'sd1810,
32'sd808, 32'sd1492, 32'sd376, 32'sd341, 32'sd630, 32'sd633,
32'sd569, 32'sd230, 32'sd1386, 32'sd1548, 32'sd325, 32'sd308,
32'sd838, 32'sd641, 32'sd1068, 32'sd148, 32'sd104, 32'sd706,
32'sd373, 32'sd247, 32'sd1875, 32'sd1649, 32'sd1486, 32'sd1135,
32'sd898, 32'sd1701, 32'sd1050, 32'sd1498, 32'sd628, 32'sd742,
32'sd1526, 32'sd435, 32'sd1331, 32'sd1066, 32'sd253, 32'sd812,
32'sd1729, 32'sd1195, 32'sd1078, 32'sd625, 32'sd225, 32'sd592,
32'sd552, 32'sd840, 32'sd479, 32'sd1284, 32'sd520, 32'sd1979,
32'sd1387, 32'sd1331, 32'sd1025, 32'sd380, 32'sd707, 32'sd1912,
32'sd1424, 32'sd1150, 32'sd1499, 32'sd1826, 32'sd547, 32'sd574,
32'sd266, 32'sd1612, 32'sd670, 32'sd817, 32'sd727, 32'sd1038,
32'sd1076, 32'sd117, 32'sd1167, 32'sd1341, 32'sd1118, 32'sd600,
32'sd1765, 32'sd1026, 32'sd979, 32'sd106, 32'sd218, 32'sd1672,
32'sd256, 32'sd1372, 32'sd291, 32'sd1771, 32'sd822, 32'sd1084,
32'sd356, 32'sd1069, 32'sd1844, 32'sd624, 32'sd1923, 32'sd1066,
32'sd1441, 32'sd713, 32'sd907, 32'sd722, 32'sd1007, 32'sd1136,
32'sd505, 32'sd1395, 32'sd1624, 32'sd517, 32'sd1855, 32'sd414,
32'sd1033, 32'sd1497, 32'sd187, 32'sd705, 32'sd1292, 32'sd283,
32'sd1553, 32'sd203, 32'sd1611, 32'sd1798, 32'sd100, 32'sd711,
32'sd1733, 32'sd1372, 32'sd1553, 32'sd1320, 32'sd1932, 32'sd693,
32'sd713, 32'sd366, 32'sd1009, 32'sd1436, 32'sd1054, 32'sd1967,
32'sd1325, 32'sd1365, 32'sd1624, 32'sd1391, 32'sd246, 32'sd1933,
32'sd458, 32'sd1690, 32'sd550, 32'sd327, 32'sd1096, 32'sd556,
32'sd1287, 32'sd705, 32'sd1485, 32'sd116, 32'sd130, 32'sd1791,
32'sd829, 32'sd183, 32'sd1344, 32'sd945, 32'sd1673, 32'sd1584,
32'sd1555, 32'sd1330, 32'sd1342, 32'sd1835, 32'sd1960, 32'sd822,
32'sd1964, 32'sd742, 32'sd999, 32'sd1788, 32'sd1276, 32'sd1969,
32'sd1966, 32'sd635, 32'sd866, 32'sd500, 32'sd1404, 32'sd832,
32'sd1919, 32'sd1044, 32'sd1064, 32'sd1336, 32'sd289, 32'sd114,
32'sd1215, 32'sd1114, 32'sd1358, 32'sd1366, 32'sd1978, 32'sd770,
32'sd1588, 32'sd642, 32'sd924, 32'sd1395, 32'sd866, 32'sd1467,
32'sd1781, 32'sd1424, 32'sd1833, 32'sd1080, 32'sd1814, 32'sd336,
32'sd374, 32'sd627, 32'sd994, 32'sd308, 32'sd1183, 32'sd725,
32'sd1968, 32'sd721, 32'sd469, 32'sd637, 32'sd1953, 32'sd885,
32'sd1630, 32'sd674, 32'sd1843, 32'sd876, 32'sd731, 32'sd1588,
32'sd249, 32'sd1649, 32'sd700, 32'sd1661, 32'sd368, 32'sd238,
32'sd534, 32'sd1532, 32'sd923, 32'sd276, 32'sd257, 32'sd1821,
32'sd1105, 32'sd1248, 32'sd787, 32'sd692, 32'sd642, 32'sd770,
32'sd1414, 32'sd1744, 32'sd886, 32'sd563, 32'sd610, 32'sd194,
32'sd883, 32'sd1461, 32'sd634, 32'sd806, 32'sd659, 32'sd1259,
32'sd126, 32'sd775, 32'sd1196, 32'sd1711, 32'sd306, 32'sd1335,
32'sd103, 32'sd1867, 32'sd936, 32'sd907, 32'sd1448, 32'sd1863,
32'sd1805, 32'sd703, 32'sd844, 32'sd1295, 32'sd277, 32'sd1910,
32'sd1488, 32'sd1297, 32'sd561, 32'sd1028, 32'sd1658, 32'sd171,
32'sd996, 32'sd1401, 32'sd759, 32'sd789, 32'sd1841, 32'sd1973,
32'sd784, 32'sd1556, 32'sd980, 32'sd681, 32'sd1177, 32'sd1267,
32'sd359, 32'sd341, 32'sd832, 32'sd1488, 32'sd1718, 32'sd1167,
32'sd1687, 32'sd583, 32'sd1522, 32'sd1434, 32'sd630, 32'sd1299,
32'sd1553, 32'sd905, 32'sd613, 32'sd938, 32'sd898, 32'sd1339,
32'sd461, 32'sd633, 32'sd1342, 32'sd1745, 32'sd1491, 32'sd133,
32'sd921, 32'sd1580, 32'sd1995, 32'sd1244, 32'sd707, 32'sd887,
32'sd1012, 32'sd622, 32'sd1589, 32'sd724, 32'sd1772, 32'sd1740,
32'sd1220, 32'sd1177, 32'sd1498, 32'sd584, 32'sd1054, 32'sd1496,
32'sd322, 32'sd1628, 32'sd446, 32'sd1630, 32'sd316, 32'sd1425,
32'sd798, 32'sd731, 32'sd1415, 32'sd1933, 32'sd1492, 32'sd1097,
32'sd1870, 32'sd1336, 32'sd981, 32'sd560, 32'sd1480, 32'sd811,
32'sd1734, 32'sd277, 32'sd290, 32'sd1969, 32'sd1469, 32'sd723,
32'sd711, 32'sd611, 32'sd252, 32'sd1882, 32'sd1877, 32'sd266,
32'sd644, 32'sd112, 32'sd925, 32'sd1275, 32'sd962, 32'sd1748,
32'sd300, 32'sd1850, 32'sd1500, 32'sd1482, 32'sd593, 32'sd522,
32'sd304, 32'sd1528, 32'sd646, 32'sd790, 32'sd1258, 32'sd1374,
32'sd708, 32'sd924, 32'sd1945, 32'sd1412, 32'sd221, 32'sd1197,
32'sd1734, 32'sd1713, 32'sd924, 32'sd1183, 32'sd862, 32'sd115,
32'sd1681, 32'sd528, 32'sd1920, 32'sd1941, 32'sd1936, 32'sd599,
32'sd322, 32'sd598, 32'sd514, 32'sd1007, 32'sd1919, 32'sd1075,
32'sd1198, 32'sd2000, 32'sd1129, 32'sd1378, 32'sd1968, 32'sd552,
32'sd211, 32'sd1219, 32'sd185, 32'sd1268, 32'sd1843, 32'sd1670,
32'sd1535, 32'sd1063, 32'sd1804, 32'sd996, 32'sd632, 32'sd421,
32'sd558, 32'sd923, 32'sd1572, 32'sd1020, 32'sd759, 32'sd103,
32'sd544, 32'sd843, 32'sd297, 32'sd1658, 32'sd876, 32'sd1361,
32'sd1404, 32'sd1514, 32'sd1483, 32'sd1275, 32'sd636, 32'sd854,
32'sd1453, 32'sd535, 32'sd1788, 32'sd898, 32'sd1136, 32'sd1212,
32'sd798, 32'sd894, 32'sd258, 32'sd643, 32'sd1660, 32'sd250,
32'sd205, 32'sd1817, 32'sd1507, 32'sd953, 32'sd1520, 32'sd1917,
32'sd1238, 32'sd574, 32'sd1148, 32'sd1226, 32'sd595, 32'sd1666,
32'sd1132, 32'sd1669, 32'sd1257, 32'sd1321, 32'sd1085, 32'sd691,
32'sd1834, 32'sd210, 32'sd149, 32'sd1375, 32'sd1911, 32'sd1532,
32'sd970, 32'sd1504, 32'sd1040, 32'sd1982, 32'sd1117, 32'sd1879,
32'sd214, 32'sd1426, 32'sd473, 32'sd1447, 32'sd1139, 32'sd297,
32'sd206, 32'sd1712, 32'sd416, 32'sd797, 32'sd1739, 32'sd1159,
32'sd1040, 32'sd112, 32'sd719, 32'sd909, 32'sd1182, 32'sd1729,
32'sd303, 32'sd622, 32'sd856, 32'sd1027, 32'sd1493, 32'sd187,
32'sd585, 32'sd347, 32'sd961, 32'sd464, 32'sd549, 32'sd1234,
32'sd666, 32'sd1874, 32'sd188, 32'sd264, 32'sd1049, 32'sd1827,
32'sd1142, 32'sd1966, 32'sd616, 32'sd1618, 32'sd335, 32'sd177,
32'sd860, 32'sd167, 32'sd1609, 32'sd248, 32'sd1638, 32'sd1380,
32'sd735, 32'sd155, 32'sd596, 32'sd544, 32'sd1463, 32'sd691,
32'sd1727, 32'sd940, 32'sd1738, 32'sd590, 32'sd791, 32'sd1450,
32'sd1950, 32'sd1551, 32'sd395, 32'sd998, 32'sd157, 32'sd1853,
32'sd800, 32'sd179, 32'sd871, 32'sd929, 32'sd1746, 32'sd1144,
32'sd1393, 32'sd1480, 32'sd1896, 32'sd520, 32'sd528, 32'sd1398,
32'sd807, 32'sd1361, 32'sd1452, 32'sd794, 32'sd1083, 32'sd814,
32'sd1606, 32'sd1765, 32'sd419, 32'sd1023, 32'sd443, 32'sd853,
32'sd1036, 32'sd1941, 32'sd1089, 32'sd147, 32'sd1171, 32'sd1398,
32'sd1258, 32'sd461, 32'sd1193, 32'sd1619, 32'sd1537, 32'sd214,
32'sd957, 32'sd1274, 32'sd1752, 32'sd1578, 32'sd498, 32'sd640,
32'sd363, 32'sd1136, 32'sd1281, 32'sd737, 32'sd1682, 32'sd1447,
32'sd1913, 32'sd1792, 32'sd1856, 32'sd1889, 32'sd697, 32'sd687,
32'sd891, 32'sd155, 32'sd1693, 32'sd100, 32'sd1404, 32'sd529,
32'sd184, 32'sd1749, 32'sd486, 32'sd827, 32'sd1278, 32'sd595,
32'sd615, 32'sd162, 32'sd1447, 32'sd685, 32'sd294, 32'sd445,
32'sd340, 32'sd1667, 32'sd1134, 32'sd230, 32'sd236, 32'sd1531,
32'sd1096, 32'sd869, 32'sd220, 32'sd881, 32'sd1024, 32'sd1829,
32'sd1546, 32'sd1661, 32'sd687, 32'sd1478, 32'sd606, 32'sd1382,
32'sd531, 32'sd1381, 32'sd1784, 32'sd1332, 32'sd922, 32'sd1667,
32'sd326, 32'sd1474, 32'sd1827, 32'sd1880, 32'sd799, 32'sd459,
32'sd684, 32'sd1166, 32'sd1974, 32'sd1351, 32'sd830, 32'sd724,
32'sd1193, 32'sd1740, 32'sd1763, 32'sd1980, 32'sd582, 32'sd825,
32'sd1907, 32'sd411, 32'sd1967, 32'sd1078, 32'sd1281, 32'sd1257,
32'sd466, 32'sd542, 32'sd756, 32'sd1690, 32'sd1420, 32'sd1723,
32'sd1752, 32'sd1640, 32'sd1069, 32'sd154, 32'sd1974, 32'sd774,
32'sd1259, 32'sd1953, 32'sd307, 32'sd194, 32'sd1283, 32'sd493,
32'sd948, 32'sd985, 32'sd127, 32'sd1243, 32'sd1750, 32'sd1412,
32'sd1437, 32'sd1440, 32'sd719, 32'sd1794, 32'sd1199, 32'sd1168,
32'sd1298, 32'sd1440, 32'sd882, 32'sd818, 32'sd1855, 32'sd510,
32'sd1567, 32'sd1320, 32'sd1018, 32'sd1632, 32'sd296, 32'sd1567,
32'sd436, 32'sd584, 32'sd1692, 32'sd990, 32'sd698, 32'sd160,
32'sd283, 32'sd1068, 32'sd180, 32'sd555, 32'sd688, 32'sd814,
32'sd267, 32'sd224, 32'sd1341, 32'sd1210, 32'sd1321, 32'sd1687,
32'sd114, 32'sd1901, 32'sd1572, 32'sd1311, 32'sd1094, 32'sd1182,
32'sd962, 32'sd1113, 32'sd1386, 32'sd1854, 32'sd857, 32'sd126,
32'sd1936, 32'sd1224, 32'sd1226, 32'sd526, 32'sd169, 32'sd1056,
32'sd595, 32'sd1243, 32'sd731, 32'sd1780, 32'sd1242, 32'sd1072,
32'sd1364, 32'sd1066, 32'sd1316, 32'sd605, 32'sd1920, 32'sd662,
32'sd627, 32'sd1570, 32'sd645, 32'sd431, 32'sd666, 32'sd157,
32'sd1739, 32'sd1570, 32'sd1271, 32'sd1083, 32'sd390, 32'sd1807,
32'sd478, 32'sd1227, 32'sd1566, 32'sd412, 32'sd1184, 32'sd514,
32'sd646, 32'sd371, 32'sd1246, 32'sd390, 32'sd1703, 32'sd381,
32'sd1854, 32'sd1506, 32'sd1692, 32'sd112, 32'sd1693, 32'sd1723,
32'sd865, 32'sd901, 32'sd552, 32'sd1341, 32'sd1643, 32'sd140,
32'sd1889, 32'sd167, 32'sd217, 32'sd857, 32'sd685, 32'sd1567,
32'sd1671, 32'sd605, 32'sd154, 32'sd1828, 32'sd1760, 32'sd1877,
32'sd1375, 32'sd1889, 32'sd561, 32'sd1363, 32'sd802, 32'sd466,
32'sd539, 32'sd142, 32'sd1806, 32'sd1632, 32'sd1086, 32'sd1653,
32'sd336, 32'sd1590, 32'sd553, 32'sd271, 32'sd899, 32'sd419,
32'sd1908, 32'sd1053, 32'sd1699, 32'sd1040, 32'sd1852, 32'sd891,
32'sd1498, 32'sd1029, 32'sd1245, 32'sd992, 32'sd411, 32'sd244,
32'sd284, 32'sd321, 32'sd1751, 32'sd1665, 32'sd1643, 32'sd288,
32'sd117, 32'sd1988, 32'sd159, 32'sd301, 32'sd1711, 32'sd1922,
32'sd490, 32'sd1403, 32'sd103, 32'sd1709, 32'sd1112, 32'sd666,
32'sd1597, 32'sd569, 32'sd999, 32'sd1966, 32'sd167, 32'sd304,
32'sd1467, 32'sd1650, 32'sd1958, 32'sd903, 32'sd1266, 32'sd1296,
32'sd398, 32'sd318, 32'sd1473, 32'sd595, 32'sd1422, 32'sd1207,
32'sd131, 32'sd1532, 32'sd1781, 32'sd1483, 32'sd1050, 32'sd924,
32'sd1787, 32'sd1076, 32'sd362, 32'sd689, 32'sd1233, 32'sd1456,
32'sd585, 32'sd1249, 32'sd1381, 32'sd1876, 32'sd1547, 32'sd1594,
32'sd1535, 32'sd1988, 32'sd525, 32'sd1431, 32'sd371, 32'sd1600,
32'sd938, 32'sd1056, 32'sd505, 32'sd1442, 32'sd1788, 32'sd1085,
32'sd1046, 32'sd354, 32'sd568, 32'sd1142, 32'sd1382, 32'sd255,
32'sd971, 32'sd1702, 32'sd985, 32'sd1091, 32'sd971, 32'sd528,
32'sd1134, 32'sd1149, 32'sd1174, 32'sd1915, 32'sd1422, 32'sd670,
32'sd784, 32'sd1601, 32'sd321, 32'sd797, 32'sd339, 32'sd176,
32'sd1075, 32'sd1049, 32'sd1035, 32'sd1256, 32'sd189, 32'sd792,
32'sd559, 32'sd1570, 32'sd352, 32'sd1339, 32'sd1485, 32'sd857,
32'sd421, 32'sd927, 32'sd1973, 32'sd1759, 32'sd1667, 32'sd1723,
32'sd555, 32'sd508, 32'sd1458, 32'sd1938, 32'sd1437, 32'sd312,
32'sd1434, 32'sd1118, 32'sd1592, 32'sd202, 32'sd816, 32'sd873,
32'sd1363, 32'sd345, 32'sd316, 32'sd1454, 32'sd1000, 32'sd731,
32'sd1666, 32'sd1761, 32'sd858, 32'sd1938, 32'sd1784, 32'sd678,
32'sd284, 32'sd446, 32'sd1270, 32'sd1031, 32'sd1058, 32'sd1635,
32'sd1172, 32'sd1209, 32'sd1166, 32'sd1392, 32'sd1976, 32'sd335,
32'sd1808, 32'sd891, 32'sd1754, 32'sd576, 32'sd1346, 32'sd1813,
32'sd1679, 32'sd1989, 32'sd1644, 32'sd1994, 32'sd440, 32'sd909,
32'sd699, 32'sd1450, 32'sd1192, 32'sd1071, 32'sd386, 32'sd1425,
32'sd1335, 32'sd448, 32'sd532, 32'sd568, 32'sd560, 32'sd438,
32'sd1413, 32'sd1768, 32'sd447, 32'sd370, 32'sd143, 32'sd1935,
32'sd485, 32'sd828, 32'sd745, 32'sd795, 32'sd451, 32'sd664,
32'sd1872, 32'sd221, 32'sd1258, 32'sd1601, 32'sd1843, 32'sd673,
32'sd950, 32'sd1053, 32'sd1698, 32'sd263, 32'sd537, 32'sd189,
32'sd844, 32'sd221, 32'sd663, 32'sd990, 32'sd651, 32'sd701,
32'sd1999, 32'sd1334, 32'sd482, 32'sd767, 32'sd297, 32'sd655,
32'sd709, 32'sd157, 32'sd1424, 32'sd1896, 32'sd298, 32'sd163,
32'sd1911, 32'sd759, 32'sd1287, 32'sd1923, 32'sd592, 32'sd981,
32'sd647, 32'sd145, 32'sd1275, 32'sd1723, 32'sd1072, 32'sd1878,
32'sd880, 32'sd1237, 32'sd990, 32'sd1864, 32'sd153, 32'sd1914,
32'sd308, 32'sd908, 32'sd511, 32'sd782, 32'sd114, 32'sd205,
32'sd1154, 32'sd270, 32'sd1385, 32'sd365, 32'sd1729, 32'sd1307,
32'sd1155, 32'sd1424, 32'sd1445, 32'sd1423, 32'sd1552, 32'sd1382,
32'sd1361, 32'sd355, 32'sd1963, 32'sd991, 32'sd1634, 32'sd1767,
32'sd131, 32'sd1120, 32'sd120, 32'sd1941, 32'sd1141, 32'sd1847,
32'sd576, 32'sd187, 32'sd541, 32'sd1176, 32'sd506, 32'sd1130,
32'sd304, 32'sd1257, 32'sd1047, 32'sd1686, 32'sd1190, 32'sd597,
32'sd1677, 32'sd888, 32'sd1518, 32'sd643, 32'sd1220, 32'sd944,
32'sd1459, 32'sd416, 32'sd1854, 32'sd1918, 32'sd1848, 32'sd1411,
32'sd1826, 32'sd1230, 32'sd948, 32'sd1494, 32'sd621, 32'sd300,
32'sd815, 32'sd832, 32'sd556, 32'sd500, 32'sd591, 32'sd356,
32'sd1593, 32'sd378, 32'sd1076, 32'sd1702, 32'sd1945, 32'sd833,
32'sd408, 32'sd472, 32'sd341, 32'sd508, 32'sd1657, 32'sd451,
32'sd668, 32'sd1244, 32'sd1006, 32'sd1649, 32'sd1061, 32'sd1272,
32'sd1460, 32'sd1059, 32'sd966, 32'sd1716, 32'sd1263, 32'sd995,
32'sd889, 32'sd1351, 32'sd1651, 32'sd483, 32'sd808, 32'sd1680,
32'sd1400, 32'sd997, 32'sd1293, 32'sd1713, 32'sd1816, 32'sd453,
32'sd249, 32'sd1824, 32'sd1771, 32'sd1239, 32'sd333, 32'sd1341,
32'sd1992, 32'sd702, 32'sd1445, 32'sd1146, 32'sd1324, 32'sd1587,
32'sd1246, 32'sd1725, 32'sd520, 32'sd468, 32'sd1074, 32'sd1943,
32'sd1233, 32'sd504, 32'sd1471, 32'sd104, 32'sd1184, 32'sd839,
32'sd577, 32'sd1427, 32'sd1117, 32'sd1883, 32'sd1061, 32'sd174,
32'sd1784, 32'sd1280, 32'sd493, 32'sd813, 32'sd1780, 32'sd1421,
32'sd1101, 32'sd890, 32'sd1669, 32'sd1552, 32'sd1609, 32'sd351,
32'sd1762, 32'sd785, 32'sd1910, 32'sd758, 32'sd1735, 32'sd1012,
32'sd1911, 32'sd1030, 32'sd1429, 32'sd1101, 32'sd1552, 32'sd1242,
32'sd1638, 32'sd1026, 32'sd1563, 32'sd1474, 32'sd1677, 32'sd1339,
32'sd1944, 32'sd1745, 32'sd377, 32'sd964, 32'sd1509, 32'sd1245,
32'sd1545, 32'sd1818, 32'sd1699, 32'sd155, 32'sd1524, 32'sd1993,
32'sd220, 32'sd213, 32'sd1731, 32'sd565, 32'sd622, 32'sd918,
32'sd1665, 32'sd1199, 32'sd692, 32'sd479, 32'sd680, 32'sd1573,
32'sd1787, 32'sd359, 32'sd1829, 32'sd281, 32'sd1610, 32'sd476,
32'sd883, 32'sd1552, 32'sd122, 32'sd460, 32'sd1609, 32'sd387,
32'sd408, 32'sd1848, 32'sd206, 32'sd1263, 32'sd1671, 32'sd459,
32'sd1908, 32'sd1211, 32'sd1942, 32'sd1130, 32'sd1160, 32'sd1451,
32'sd928, 32'sd384, 32'sd1902, 32'sd1407, 32'sd796, 32'sd1636,
32'sd1285, 32'sd485, 32'sd713, 32'sd1716, 32'sd845, 32'sd1855,
32'sd1564, 32'sd1380, 32'sd984, 32'sd1967, 32'sd1004, 32'sd1282,
32'sd1931, 32'sd1997, 32'sd473, 32'sd353, 32'sd1494, 32'sd262,
32'sd1185, 32'sd333, 32'sd1462, 32'sd1775, 32'sd1868, 32'sd1684,
32'sd1025, 32'sd874, 32'sd1810, 32'sd1023, 32'sd380, 32'sd607,
32'sd1715, 32'sd1808, 32'sd219, 32'sd245, 32'sd1561, 32'sd1014,
32'sd360, 32'sd1698, 32'sd1328, 32'sd1356, 32'sd776, 32'sd504,
32'sd442, 32'sd382, 32'sd231, 32'sd992, 32'sd1813, 32'sd103,
32'sd643, 32'sd1037, 32'sd217, 32'sd1278, 32'sd1285, 32'sd598,
32'sd1821, 32'sd1965, 32'sd315, 32'sd1241, 32'sd1680, 32'sd1465,
32'sd243, 32'sd1940, 32'sd1771, 32'sd2000, 32'sd574, 32'sd1030,
32'sd1690, 32'sd1661, 32'sd1459, 32'sd1593, 32'sd930, 32'sd1209,
32'sd502, 32'sd649, 32'sd233, 32'sd197, 32'sd1636, 32'sd790,
32'sd1678, 32'sd1023, 32'sd349, 32'sd409, 32'sd1060, 32'sd532,
32'sd633, 32'sd1572, 32'sd1419, 32'sd1515, 32'sd1975, 32'sd1225,
32'sd1320, 32'sd269, 32'sd1565, 32'sd1330, 32'sd829, 32'sd723,
32'sd256, 32'sd733, 32'sd1760, 32'sd1830, 32'sd1467, 32'sd1593,
32'sd1895, 32'sd1344, 32'sd1977, 32'sd186, 32'sd1467, 32'sd1268,
32'sd951, 32'sd1816, 32'sd562, 32'sd1654, 32'sd1467, 32'sd1780,
32'sd1472, 32'sd1558, 32'sd271, 32'sd1593, 32'sd1923, 32'sd1329,
32'sd1467, 32'sd228, 32'sd739, 32'sd790, 32'sd578, 32'sd539,
32'sd1903, 32'sd1361, 32'sd285, 32'sd1109, 32'sd1812, 32'sd1633,
32'sd1011, 32'sd827, 32'sd1983, 32'sd1134, 32'sd674, 32'sd226,
32'sd1220, 32'sd1162, 32'sd1308, 32'sd681, 32'sd1533, 32'sd1952,
32'sd726, 32'sd747, 32'sd674, 32'sd1860, 32'sd1683, 32'sd1270,
32'sd1729, 32'sd1964, 32'sd1428, 32'sd536, 32'sd1178, 32'sd358,
32'sd1284, 32'sd1176, 32'sd638, 32'sd1195, 32'sd1063, 32'sd1696,
32'sd1496, 32'sd1898, 32'sd1149, 32'sd1157, 32'sd1907, 32'sd785,
32'sd634, 32'sd1379, 32'sd290, 32'sd1870, 32'sd1646, 32'sd148,
32'sd104, 32'sd1344, 32'sd479, 32'sd815, 32'sd1812, 32'sd428,
32'sd419, 32'sd1129, 32'sd707, 32'sd1305, 32'sd1657, 32'sd967,
32'sd1089, 32'sd635, 32'sd1276, 32'sd749, 32'sd1538, 32'sd1952,
32'sd364, 32'sd1158, 32'sd1589, 32'sd1760, 32'sd799, 32'sd819,
32'sd146, 32'sd1568, 32'sd841, 32'sd543, 32'sd670, 32'sd746,
32'sd1019, 32'sd273, 32'sd389, 32'sd1149, 32'sd147, 32'sd106,
32'sd730, 32'sd802, 32'sd1288, 32'sd1520, 32'sd1679, 32'sd1622,
32'sd1764, 32'sd1502, 32'sd643, 32'sd517, 32'sd1619, 32'sd684,
32'sd760, 32'sd471, 32'sd1510, 32'sd1838, 32'sd1709, 32'sd621,
32'sd1975, 32'sd312, 32'sd985, 32'sd405, 32'sd421, 32'sd1353,
32'sd1382, 32'sd1184, 32'sd173, 32'sd206, 32'sd558, 32'sd1229,
32'sd1233, 32'sd1028, 32'sd1418, 32'sd1140, 32'sd1797, 32'sd259,
32'sd1993, 32'sd748, 32'sd1863, 32'sd1916, 32'sd956, 32'sd635,
32'sd375, 32'sd974, 32'sd559, 32'sd870, 32'sd820, 32'sd1786,
32'sd586, 32'sd448, 32'sd866, 32'sd1547, 32'sd1053, 32'sd778,
32'sd102, 32'sd1683, 32'sd921, 32'sd1336, 32'sd124, 32'sd475,
32'sd569, 32'sd416, 32'sd187, 32'sd1264, 32'sd244, 32'sd571,
32'sd436, 32'sd1586, 32'sd1673, 32'sd1826, 32'sd491, 32'sd1432,
32'sd443, 32'sd1574, 32'sd398, 32'sd238, 32'sd1620, 32'sd351,
32'sd1266, 32'sd1782, 32'sd703, 32'sd1250, 32'sd1615, 32'sd983,
32'sd1553, 32'sd565, 32'sd916, 32'sd1655, 32'sd1240, 32'sd570,
32'sd1481, 32'sd583, 32'sd189, 32'sd234, 32'sd743, 32'sd1063,
32'sd1860, 32'sd1805, 32'sd1765, 32'sd1376, 32'sd1002, 32'sd1275,
32'sd1828, 32'sd658, 32'sd658, 32'sd580, 32'sd1969, 32'sd1748,
32'sd640, 32'sd836, 32'sd263, 32'sd541, 32'sd192, 32'sd1734,
32'sd1836, 32'sd977, 32'sd990, 32'sd521, 32'sd1960, 32'sd803,
32'sd781, 32'sd927, 32'sd971, 32'sd1771, 32'sd157, 32'sd729,
32'sd1163, 32'sd134, 32'sd1526, 32'sd962, 32'sd626, 32'sd1892,
32'sd1282, 32'sd220, 32'sd199, 32'sd900, 32'sd1630, 32'sd1455,
32'sd1116, 32'sd1845, 32'sd536, 32'sd698, 32'sd1378, 32'sd1147,
32'sd499, 32'sd725, 32'sd1654, 32'sd1433, 32'sd992, 32'sd244,
32'sd1257, 32'sd1355, 32'sd415, 32'sd1180, 32'sd465, 32'sd1260,
32'sd537, 32'sd1034, 32'sd854, 32'sd1708, 32'sd1473, 32'sd1417,
32'sd432, 32'sd1357, 32'sd813, 32'sd618, 32'sd562, 32'sd1174,
32'sd116, 32'sd524, 32'sd1720, 32'sd1496, 32'sd1368, 32'sd537,
32'sd1598, 32'sd1402, 32'sd247, 32'sd1540, 32'sd1527, 32'sd1472,
32'sd1617, 32'sd1355, 32'sd943, 32'sd412, 32'sd278, 32'sd1653,
32'sd539, 32'sd459, 32'sd536, 32'sd1005, 32'sd1216, 32'sd1305,
32'sd1505, 32'sd1208, 32'sd1060, 32'sd956, 32'sd1242, 32'sd1745,
32'sd110, 32'sd1634, 32'sd1561, 32'sd768, 32'sd1358, 32'sd1846,
32'sd348, 32'sd1295, 32'sd753, 32'sd1028, 32'sd783, 32'sd245,
32'sd872, 32'sd1301, 32'sd569, 32'sd1629, 32'sd1357, 32'sd684,
32'sd315, 32'sd321, 32'sd514, 32'sd783, 32'sd1622, 32'sd846,
32'sd1359, 32'sd1295, 32'sd224, 32'sd1025, 32'sd1244, 32'sd1927,
32'sd1110, 32'sd498, 32'sd1060, 32'sd1058, 32'sd1395, 32'sd991,
32'sd1581, 32'sd908, 32'sd1514, 32'sd1491, 32'sd1427, 32'sd125,
32'sd1708, 32'sd440, 32'sd1684, 32'sd619, 32'sd1043, 32'sd1763,
32'sd1700, 32'sd374, 32'sd565, 32'sd1613, 32'sd1998, 32'sd1084,
32'sd1773, 32'sd125, 32'sd1066, 32'sd1506, 32'sd818, 32'sd1305,
32'sd682, 32'sd1557, 32'sd252, 32'sd117, 32'sd381, 32'sd406,
32'sd512, 32'sd1988, 32'sd713, 32'sd1593, 32'sd123, 32'sd1838,
32'sd495, 32'sd278, 32'sd766, 32'sd557, 32'sd156, 32'sd902,
32'sd1043, 32'sd519, 32'sd883, 32'sd1689, 32'sd1998, 32'sd1519,
32'sd300, 32'sd1017, 32'sd1375, 32'sd1722, 32'sd163, 32'sd1071,
32'sd1929, 32'sd1041, 32'sd332, 32'sd104, 32'sd1195, 32'sd1477,
32'sd476, 32'sd1850, 32'sd533, 32'sd1280, 32'sd172, 32'sd621,
32'sd166, 32'sd1866, 32'sd152, 32'sd1164, 32'sd1530, 32'sd1125,
32'sd858, 32'sd1804, 32'sd1886, 32'sd351, 32'sd1099, 32'sd1509,
32'sd513, 32'sd1174, 32'sd527, 32'sd1661, 32'sd1456, 32'sd1431,
32'sd1517, 32'sd1403, 32'sd104, 32'sd756, 32'sd972, 32'sd1978,
32'sd830, 32'sd873, 32'sd136, 32'sd1561, 32'sd712, 32'sd877,
32'sd229, 32'sd265, 32'sd498, 32'sd901, 32'sd1099, 32'sd201,
32'sd1832, 32'sd1537, 32'sd1737, 32'sd265, 32'sd159, 32'sd958,
32'sd1315, 32'sd1412, 32'sd1714, 32'sd672, 32'sd822, 32'sd1289,
32'sd926, 32'sd409, 32'sd497, 32'sd756, 32'sd870, 32'sd1417,
32'sd266, 32'sd1495, 32'sd980, 32'sd419, 32'sd245, 32'sd1439,
32'sd707, 32'sd599, 32'sd1691, 32'sd248, 32'sd679, 32'sd1686,
32'sd706, 32'sd418, 32'sd491, 32'sd728, 32'sd1437, 32'sd338,
32'sd1767, 32'sd751, 32'sd1991, 32'sd267, 32'sd928, 32'sd367,
32'sd321, 32'sd893, 32'sd1888, 32'sd1292, 32'sd1614, 32'sd1657,
32'sd1652, 32'sd424, 32'sd926, 32'sd1766, 32'sd786, 32'sd215,
32'sd1463, 32'sd1801, 32'sd480, 32'sd920, 32'sd1587, 32'sd1142,
32'sd706, 32'sd1689, 32'sd509, 32'sd1343, 32'sd1435, 32'sd1800,
32'sd1691, 32'sd639, 32'sd1210, 32'sd461, 32'sd256, 32'sd1614,
32'sd760, 32'sd281, 32'sd281, 32'sd1287, 32'sd1226, 32'sd135,
32'sd1501, 32'sd1601, 32'sd1777, 32'sd558, 32'sd1099, 32'sd1847,
32'sd142, 32'sd511, 32'sd776, 32'sd1262, 32'sd1271, 32'sd928,
32'sd1835, 32'sd1020, 32'sd785, 32'sd200, 32'sd892, 32'sd554,
32'sd1090, 32'sd177, 32'sd1036, 32'sd229, 32'sd984, 32'sd824,
32'sd1819, 32'sd1344, 32'sd1585, 32'sd640, 32'sd1198, 32'sd1155,
32'sd194, 32'sd1834, 32'sd577, 32'sd1662, 32'sd1549, 32'sd1388,
32'sd1149, 32'sd1643, 32'sd872, 32'sd1411, 32'sd1272, 32'sd146,
32'sd422, 32'sd1902, 32'sd190, 32'sd443, 32'sd1739, 32'sd1925,
32'sd1780, 32'sd1680, 32'sd202, 32'sd1366, 32'sd1592, 32'sd1198,
32'sd1801, 32'sd1918, 32'sd303, 32'sd1285, 32'sd1478, 32'sd1175,
32'sd1688, 32'sd731, 32'sd885, 32'sd1882, 32'sd285, 32'sd945,
32'sd297, 32'sd355, 32'sd1325, 32'sd1592, 32'sd1237, 32'sd725,
32'sd1956, 32'sd1096, 32'sd1450, 32'sd133, 32'sd1730, 32'sd673,
32'sd279, 32'sd1413, 32'sd1210, 32'sd460, 32'sd223, 32'sd1373,
32'sd1097, 32'sd303, 32'sd1600, 32'sd1942, 32'sd1359, 32'sd1678,
32'sd1980, 32'sd331, 32'sd1048, 32'sd1591, 32'sd1645, 32'sd1152,
32'sd1491, 32'sd1542, 32'sd806, 32'sd988, 32'sd1329, 32'sd506,
32'sd537, 32'sd1964, 32'sd206, 32'sd167, 32'sd1807, 32'sd1608,
32'sd1297, 32'sd277, 32'sd111, 32'sd934, 32'sd222, 32'sd1187,
32'sd198, 32'sd838, 32'sd1225, 32'sd894, 32'sd1261, 32'sd752,
32'sd1520, 32'sd901, 32'sd692, 32'sd1977, 32'sd1910, 32'sd554,
32'sd772, 32'sd820, 32'sd964, 32'sd612, 32'sd488, 32'sd1764,
32'sd1129, 32'sd177, 32'sd938, 32'sd661, 32'sd946, 32'sd1991,
32'sd1235, 32'sd456, 32'sd1690, 32'sd1246, 32'sd1845, 32'sd1493,
32'sd241, 32'sd1425, 32'sd1216, 32'sd671, 32'sd1111, 32'sd110,
32'sd1679, 32'sd1104, 32'sd869, 32'sd1715, 32'sd320, 32'sd1811,
32'sd1835, 32'sd232, 32'sd1725, 32'sd135, 32'sd1888, 32'sd393,
32'sd1695, 32'sd1030, 32'sd1914, 32'sd786, 32'sd1801, 32'sd1627,
32'sd280, 32'sd453, 32'sd1796, 32'sd202, 32'sd235, 32'sd1255,
32'sd1502, 32'sd1069, 32'sd1370, 32'sd1798, 32'sd1228, 32'sd1824,
32'sd1820, 32'sd285, 32'sd1990, 32'sd1975, 32'sd272, 32'sd1968,
32'sd364, 32'sd448, 32'sd1847, 32'sd1331, 32'sd313, 32'sd1062,
32'sd1519, 32'sd1828, 32'sd1118, 32'sd1492, 32'sd1081, 32'sd1565,
32'sd250, 32'sd434, 32'sd220, 32'sd731, 32'sd1377, 32'sd949,
32'sd1269, 32'sd1242, 32'sd1956, 32'sd628, 32'sd616, 32'sd1340,
32'sd586, 32'sd262, 32'sd973, 32'sd1667, 32'sd347, 32'sd1182,
32'sd251, 32'sd933, 32'sd1913, 32'sd1820, 32'sd1479, 32'sd1164,
32'sd1844, 32'sd704, 32'sd928, 32'sd1118, 32'sd1915, 32'sd1909,
32'sd742, 32'sd787, 32'sd1121, 32'sd1550, 32'sd1837, 32'sd1572,
32'sd112, 32'sd1276, 32'sd643, 32'sd786, 32'sd1277, 32'sd228,
32'sd1499, 32'sd400, 32'sd1560, 32'sd1054, 32'sd191, 32'sd1865,
32'sd275, 32'sd881, 32'sd1042, 32'sd1824, 32'sd482, 32'sd1512,
32'sd1920, 32'sd631, 32'sd134, 32'sd368, 32'sd567, 32'sd194,
32'sd1820, 32'sd1004, 32'sd606, 32'sd1943, 32'sd120, 32'sd933,
32'sd144, 32'sd566, 32'sd428, 32'sd563, 32'sd134, 32'sd366,
32'sd532, 32'sd787, 32'sd802, 32'sd229, 32'sd701, 32'sd482,
32'sd1454, 32'sd1446, 32'sd482, 32'sd1251, 32'sd1830, 32'sd1623,
32'sd299, 32'sd1559, 32'sd852, 32'sd512, 32'sd1584, 32'sd704,
32'sd1239, 32'sd221, 32'sd295, 32'sd514, 32'sd450, 32'sd1700,
32'sd183, 32'sd1138, 32'sd1105, 32'sd124, 32'sd1810, 32'sd1579,
32'sd1954, 32'sd1672, 32'sd217, 32'sd1773, 32'sd1625, 32'sd1353,
32'sd609, 32'sd925, 32'sd1517, 32'sd563, 32'sd577, 32'sd1432,
32'sd713, 32'sd1457, 32'sd869, 32'sd823, 32'sd1232, 32'sd560,
32'sd1797, 32'sd209, 32'sd1529, 32'sd854, 32'sd669, 32'sd1725,
32'sd993, 32'sd1911, 32'sd1420, 32'sd531, 32'sd109, 32'sd1989,
32'sd1971, 32'sd343, 32'sd1085, 32'sd1022, 32'sd756, 32'sd759,
32'sd1132, 32'sd1646, 32'sd793, 32'sd893, 32'sd847, 32'sd728,
32'sd186, 32'sd1141, 32'sd917, 32'sd1854, 32'sd1607, 32'sd1567,
32'sd872, 32'sd1593, 32'sd940, 32'sd1125, 32'sd672, 32'sd1619,
32'sd129, 32'sd1818, 32'sd530, 32'sd1694, 32'sd1210, 32'sd176,
32'sd1459, 32'sd692, 32'sd1087, 32'sd1482, 32'sd144, 32'sd1785,
32'sd1904, 32'sd491, 32'sd1968, 32'sd1703, 32'sd1814, 32'sd1654,
32'sd794, 32'sd820, 32'sd663, 32'sd273, 32'sd1242, 32'sd917,
32'sd849, 32'sd1168, 32'sd1672, 32'sd844, 32'sd1770, 32'sd151,
32'sd893, 32'sd1860, 32'sd119, 32'sd485, 32'sd1305, 32'sd1654,
32'sd1986, 32'sd181, 32'sd451, 32'sd1338, 32'sd1139, 32'sd615,
32'sd1822, 32'sd1442, 32'sd1535, 32'sd196, 32'sd574, 32'sd665,
32'sd1774, 32'sd1566, 32'sd1316, 32'sd608, 32'sd1727, 32'sd514,
32'sd1914, 32'sd720, 32'sd1026, 32'sd801, 32'sd753, 32'sd856,
32'sd311, 32'sd349, 32'sd484, 32'sd1972, 32'sd405, 32'sd1496,
32'sd760, 32'sd1968, 32'sd1573, 32'sd1151, 32'sd799, 32'sd1328,
32'sd1398, 32'sd1624, 32'sd938, 32'sd1138, 32'sd173, 32'sd617,
32'sd422, 32'sd487, 32'sd535, 32'sd122, 32'sd962, 32'sd901,
32'sd1231, 32'sd1560, 32'sd1343, 32'sd968, 32'sd931, 32'sd518,
32'sd1319, 32'sd442, 32'sd1062, 32'sd1551, 32'sd338, 32'sd754,
32'sd1891, 32'sd601, 32'sd923, 32'sd1247, 32'sd175, 32'sd350,
32'sd311, 32'sd145, 32'sd185, 32'sd503, 32'sd1399, 32'sd1330,
32'sd1262, 32'sd981, 32'sd659, 32'sd1105, 32'sd719, 32'sd399,
32'sd1010, 32'sd385, 32'sd1106, 32'sd897, 32'sd809, 32'sd1310,
32'sd1317, 32'sd719, 32'sd893, 32'sd1176, 32'sd1169, 32'sd906,
32'sd1909, 32'sd986, 32'sd1082, 32'sd1877, 32'sd1482, 32'sd1478,
32'sd1483, 32'sd1488, 32'sd730, 32'sd1181, 32'sd872, 32'sd163,
32'sd1483, 32'sd447, 32'sd1876, 32'sd1689, 32'sd1001, 32'sd330,
32'sd1349, 32'sd850, 32'sd1840, 32'sd299, 32'sd1138, 32'sd416,
32'sd933, 32'sd442, 32'sd1018, 32'sd1071, 32'sd899, 32'sd1539,
32'sd1632, 32'sd1338, 32'sd1780, 32'sd1164, 32'sd920, 32'sd646,
32'sd1457, 32'sd1288, 32'sd1056, 32'sd1974, 32'sd1133, 32'sd1480,
32'sd1116, 32'sd555, 32'sd805, 32'sd790, 32'sd653, 32'sd1687,
32'sd1614, 32'sd132, 32'sd1270, 32'sd532, 32'sd1065, 32'sd519,
32'sd735, 32'sd277, 32'sd219, 32'sd1438, 32'sd1210, 32'sd860,
32'sd1789, 32'sd1296, 32'sd1082, 32'sd1774, 32'sd1025, 32'sd1376,
32'sd1170, 32'sd1014, 32'sd293, 32'sd1558, 32'sd1701, 32'sd1104,
32'sd1617, 32'sd1495, 32'sd944, 32'sd775, 32'sd1778, 32'sd898,
32'sd649, 32'sd662, 32'sd592, 32'sd386, 32'sd963, 32'sd1218,
32'sd765, 32'sd842, 32'sd1396, 32'sd942, 32'sd1676, 32'sd1149,
32'sd740, 32'sd124, 32'sd998, 32'sd1876, 32'sd1002, 32'sd1142,
32'sd1873, 32'sd1911, 32'sd225, 32'sd931, 32'sd1044, 32'sd1577,
32'sd536, 32'sd372, 32'sd632, 32'sd965, 32'sd1030, 32'sd1815,
32'sd1876, 32'sd1969, 32'sd1015, 32'sd1592, 32'sd505, 32'sd609,
32'sd1327, 32'sd1987, 32'sd1734, 32'sd460, 32'sd973, 32'sd799,
32'sd1615, 32'sd1396, 32'sd327, 32'sd1785, 32'sd517, 32'sd1305,
32'sd1994, 32'sd844, 32'sd1626, 32'sd1671, 32'sd878, 32'sd1283,
32'sd1372, 32'sd1384, 32'sd1087, 32'sd1518, 32'sd122, 32'sd468,
32'sd1539, 32'sd1433, 32'sd1380, 32'sd274, 32'sd148, 32'sd1802,
32'sd1585, 32'sd519, 32'sd212, 32'sd145, 32'sd918, 32'sd930,
32'sd1515, 32'sd1571, 32'sd462, 32'sd1213, 32'sd537, 32'sd1359,
32'sd794, 32'sd1453, 32'sd1771, 32'sd488, 32'sd1831, 32'sd1811,
32'sd1542, 32'sd1966, 32'sd1939, 32'sd498, 32'sd1242, 32'sd964,
32'sd249, 32'sd1831, 32'sd1909, 32'sd408, 32'sd734, 32'sd710,
32'sd1432, 32'sd1148, 32'sd138, 32'sd1308, 32'sd628, 32'sd567,
32'sd545, 32'sd827, 32'sd1889, 32'sd907, 32'sd1489, 32'sd1270,
32'sd463, 32'sd417, 32'sd1150, 32'sd1431, 32'sd1928, 32'sd560,
32'sd1821, 32'sd1288, 32'sd429, 32'sd668, 32'sd488, 32'sd1367,
32'sd1223, 32'sd698, 32'sd940, 32'sd1550, 32'sd508, 32'sd742,
32'sd184, 32'sd350, 32'sd120, 32'sd182, 32'sd1511, 32'sd136,
32'sd283, 32'sd1581, 32'sd865, 32'sd1213, 32'sd1559, 32'sd1555,
32'sd1801, 32'sd1512, 32'sd1377, 32'sd1200, 32'sd1567, 32'sd313,
32'sd1824, 32'sd546, 32'sd279, 32'sd253, 32'sd116, 32'sd576,
32'sd932, 32'sd1029, 32'sd1717, 32'sd1178, 32'sd1739, 32'sd1452,
32'sd743, 32'sd197, 32'sd327, 32'sd964, 32'sd1951, 32'sd651,
32'sd1462, 32'sd1245, 32'sd1783, 32'sd1295, 32'sd1027, 32'sd1352,
32'sd197, 32'sd1376, 32'sd1430, 32'sd1146, 32'sd1667, 32'sd1749,
32'sd1537, 32'sd368, 32'sd636, 32'sd1041, 32'sd647, 32'sd1494,
32'sd1586, 32'sd1803, 32'sd247, 32'sd1971, 32'sd1411, 32'sd1740,
32'sd889, 32'sd1564, 32'sd723, 32'sd493, 32'sd149, 32'sd264,
32'sd1354, 32'sd483, 32'sd732, 32'sd724, 32'sd1464, 32'sd1135,
32'sd1353, 32'sd1265, 32'sd1266, 32'sd182, 32'sd515, 32'sd1950,
32'sd433, 32'sd1528, 32'sd1097, 32'sd976, 32'sd211, 32'sd581,
32'sd1149, 32'sd1652, 32'sd1576, 32'sd1332, 32'sd1109, 32'sd369,
32'sd1634, 32'sd1501, 32'sd326, 32'sd342, 32'sd1099, 32'sd212,
32'sd550, 32'sd1065, 32'sd274, 32'sd389, 32'sd446, 32'sd990,
32'sd913, 32'sd1130, 32'sd869, 32'sd1400, 32'sd1084, 32'sd1341,
32'sd399, 32'sd1063, 32'sd222, 32'sd1412, 32'sd576, 32'sd1283,
32'sd1157, 32'sd306, 32'sd593, 32'sd707, 32'sd1481, 32'sd1936,
32'sd1530, 32'sd159, 32'sd1480, 32'sd1952, 32'sd1788, 32'sd1992,
32'sd1096, 32'sd904, 32'sd1369, 32'sd1788, 32'sd464, 32'sd238,
32'sd156, 32'sd1020, 32'sd651, 32'sd862, 32'sd916, 32'sd336,
32'sd1818, 32'sd1360, 32'sd1089, 32'sd196, 32'sd832, 32'sd1908,
32'sd112, 32'sd188, 32'sd369, 32'sd857, 32'sd1508, 32'sd298,
32'sd1540, 32'sd962, 32'sd1127, 32'sd111, 32'sd1267, 32'sd1337,
32'sd964, 32'sd935, 32'sd621, 32'sd1827, 32'sd479, 32'sd1116,
32'sd1699, 32'sd1564, 32'sd1008, 32'sd576, 32'sd649, 32'sd1233,
32'sd1454, 32'sd1052, 32'sd1743, 32'sd834, 32'sd1301, 32'sd551,
32'sd817, 32'sd653, 32'sd1239, 32'sd111, 32'sd1187, 32'sd1489,
32'sd825, 32'sd1465, 32'sd615, 32'sd838, 32'sd1706, 32'sd1454,
32'sd1774, 32'sd1346, 32'sd283, 32'sd1329, 32'sd470, 32'sd1078,
32'sd1705, 32'sd1034, 32'sd1143, 32'sd150, 32'sd304, 32'sd1903,
32'sd1771, 32'sd761, 32'sd194, 32'sd674, 32'sd380, 32'sd165,
32'sd1261, 32'sd406, 32'sd1658, 32'sd618, 32'sd406, 32'sd1153,
32'sd1638, 32'sd607, 32'sd855, 32'sd1543, 32'sd1256, 32'sd488,
32'sd306, 32'sd1975, 32'sd1324, 32'sd925, 32'sd1318, 32'sd252,
32'sd760, 32'sd163, 32'sd1973, 32'sd219, 32'sd1928, 32'sd484,
32'sd732, 32'sd1151, 32'sd543, 32'sd1928, 32'sd1492, 32'sd597,
32'sd1193, 32'sd668, 32'sd1057, 32'sd452, 32'sd853, 32'sd125,
32'sd889, 32'sd263, 32'sd140, 32'sd1676, 32'sd1808, 32'sd1980,
32'sd1090, 32'sd1007, 32'sd1144, 32'sd315, 32'sd498, 32'sd1814,
32'sd781, 32'sd724, 32'sd704, 32'sd1026, 32'sd459, 32'sd964,
32'sd299, 32'sd315, 32'sd696, 32'sd1300, 32'sd346, 32'sd267,
32'sd408, 32'sd659, 32'sd1573, 32'sd1474, 32'sd713, 32'sd1273,
32'sd415, 32'sd1366, 32'sd935, 32'sd620, 32'sd1448, 32'sd515,
32'sd1832, 32'sd1925, 32'sd169, 32'sd1684, 32'sd811, 32'sd516,
32'sd406, 32'sd1446, 32'sd1195, 32'sd584, 32'sd970, 32'sd1161,
32'sd1967, 32'sd434, 32'sd1434, 32'sd1912, 32'sd200, 32'sd1744,
32'sd1908, 32'sd615, 32'sd682, 32'sd1383, 32'sd1420, 32'sd1061,
32'sd1796, 32'sd361, 32'sd130, 32'sd690, 32'sd497, 32'sd423,
32'sd1051, 32'sd1504, 32'sd1715, 32'sd700, 32'sd592, 32'sd1388,
32'sd1810, 32'sd738, 32'sd1500, 32'sd691, 32'sd1677, 32'sd1907,
32'sd1624, 32'sd1640, 32'sd1662, 32'sd244, 32'sd1744, 32'sd795,
32'sd1303, 32'sd482, 32'sd985, 32'sd1950, 32'sd1216, 32'sd842,
32'sd1307, 32'sd589, 32'sd421, 32'sd565, 32'sd1297, 32'sd322,
32'sd1159, 32'sd378, 32'sd1617, 32'sd809, 32'sd1141, 32'sd967,
32'sd1925, 32'sd1215, 32'sd541, 32'sd1738, 32'sd324, 32'sd281,
32'sd1811, 32'sd702, 32'sd539, 32'sd1059, 32'sd147, 32'sd983,
32'sd1361, 32'sd713, 32'sd1413, 32'sd1806, 32'sd1791, 32'sd1168,
32'sd1571, 32'sd1787, 32'sd1548, 32'sd877, 32'sd450, 32'sd211,
32'sd1202, 32'sd348, 32'sd1190, 32'sd1680, 32'sd1044, 32'sd1162,
32'sd1837, 32'sd478, 32'sd1763, 32'sd1771, 32'sd1804, 32'sd1542,
32'sd657, 32'sd891, 32'sd327, 32'sd923, 32'sd734, 32'sd480,
32'sd1126, 32'sd212, 32'sd1201, 32'sd600, 32'sd451, 32'sd1737,
32'sd1710, 32'sd849, 32'sd1617, 32'sd1349, 32'sd406, 32'sd1212,
32'sd1200, 32'sd183, 32'sd424, 32'sd1422, 32'sd1674, 32'sd861,
32'sd1075, 32'sd1753, 32'sd247, 32'sd1832, 32'sd1741, 32'sd1439,
32'sd894, 32'sd706, 32'sd1012, 32'sd1461, 32'sd393, 32'sd1642,
32'sd837, 32'sd1455, 32'sd528, 32'sd434, 32'sd837, 32'sd1848,
32'sd136, 32'sd1876, 32'sd1314, 32'sd1566, 32'sd1554, 32'sd462,
32'sd693, 32'sd992, 32'sd1196, 32'sd1733, 32'sd1215, 32'sd1545,
32'sd1208, 32'sd580, 32'sd1886, 32'sd313, 32'sd582, 32'sd1888,
32'sd1978, 32'sd1442, 32'sd180, 32'sd1974, 32'sd372, 32'sd1960,
32'sd418, 32'sd841, 32'sd1416, 32'sd468, 32'sd1179, 32'sd1155,
32'sd526, 32'sd840, 32'sd169, 32'sd1638, 32'sd1950, 32'sd1613,
32'sd1058, 32'sd789, 32'sd972, 32'sd1223, 32'sd1439, 32'sd822,
32'sd1337, 32'sd695, 32'sd1528, 32'sd1314, 32'sd454, 32'sd200,
32'sd1259, 32'sd1557, 32'sd646, 32'sd1105, 32'sd1424, 32'sd1775,
32'sd266, 32'sd750, 32'sd344, 32'sd871, 32'sd1294, 32'sd945,
32'sd1110, 32'sd1572, 32'sd329, 32'sd1153, 32'sd1309, 32'sd1602,
32'sd1860, 32'sd1184, 32'sd251, 32'sd312, 32'sd260, 32'sd1696,
32'sd285, 32'sd409, 32'sd1850, 32'sd814, 32'sd897, 32'sd392,
32'sd1715, 32'sd383, 32'sd1948, 32'sd1866, 32'sd713, 32'sd1560,
32'sd1516, 32'sd1216, 32'sd892, 32'sd1528, 32'sd150, 32'sd1691,
32'sd1518, 32'sd812, 32'sd343, 32'sd1665, 32'sd1233, 32'sd1961,
32'sd1602, 32'sd1134, 32'sd1862, 32'sd1743, 32'sd939, 32'sd895,
32'sd1103, 32'sd624, 32'sd376, 32'sd268, 32'sd281, 32'sd316,
32'sd1081, 32'sd1580, 32'sd1938, 32'sd1771, 32'sd266, 32'sd1592,
32'sd1512, 32'sd627, 32'sd1683, 32'sd1666, 32'sd946, 32'sd986,
32'sd521, 32'sd1697, 32'sd1261, 32'sd1453, 32'sd1348, 32'sd1623,
32'sd1053, 32'sd1275, 32'sd1284, 32'sd190, 32'sd110, 32'sd1737,
32'sd861, 32'sd1864, 32'sd727, 32'sd619, 32'sd405, 32'sd658,
32'sd1779, 32'sd284, 32'sd673, 32'sd686, 32'sd734, 32'sd659,
32'sd841, 32'sd1285, 32'sd703, 32'sd1813, 32'sd1460, 32'sd741,
32'sd1026, 32'sd854, 32'sd1983, 32'sd381, 32'sd1052, 32'sd203,
32'sd775, 32'sd1373, 32'sd289, 32'sd141, 32'sd1583, 32'sd418,
32'sd262, 32'sd1595, 32'sd346, 32'sd1321, 32'sd159, 32'sd622,
32'sd1355, 32'sd363, 32'sd1735, 32'sd169, 32'sd1893, 32'sd1023,
32'sd1340, 32'sd103, 32'sd874, 32'sd1917, 32'sd671, 32'sd648,
32'sd1949, 32'sd1618, 32'sd1373, 32'sd1305, 32'sd604, 32'sd1940,
32'sd349, 32'sd723, 32'sd843, 32'sd1736, 32'sd1612, 32'sd1530,
32'sd1345, 32'sd1712, 32'sd1089, 32'sd1583, 32'sd1472, 32'sd626,
32'sd387, 32'sd1226, 32'sd1964, 32'sd575, 32'sd1290, 32'sd1295,
32'sd1346, 32'sd1972, 32'sd1293, 32'sd347, 32'sd1531, 32'sd1215,
32'sd716, 32'sd713, 32'sd879, 32'sd1797, 32'sd1350, 32'sd1841,
32'sd1510, 32'sd1467, 32'sd1395, 32'sd1643, 32'sd365, 32'sd375,
32'sd241, 32'sd730, 32'sd604, 32'sd1783, 32'sd1376, 32'sd835,
32'sd1997, 32'sd1141, 32'sd627, 32'sd1967, 32'sd578, 32'sd197,
32'sd1863, 32'sd318, 32'sd1777, 32'sd288, 32'sd1678, 32'sd853,
32'sd1110, 32'sd1672, 32'sd1959, 32'sd102, 32'sd821, 32'sd1388,
32'sd1506, 32'sd1071, 32'sd363, 32'sd454, 32'sd1397, 32'sd348,
32'sd1691, 32'sd966, 32'sd869, 32'sd1831, 32'sd1996, 32'sd1878,
32'sd143, 32'sd684, 32'sd854, 32'sd1109, 32'sd503, 32'sd570,
32'sd207, 32'sd1824, 32'sd817, 32'sd1634, 32'sd154, 32'sd493,
32'sd1402, 32'sd1841, 32'sd1540, 32'sd1138, 32'sd1474, 32'sd742,
32'sd1421, 32'sd343, 32'sd815, 32'sd463, 32'sd467, 32'sd432,
32'sd786, 32'sd1099, 32'sd1074, 32'sd856, 32'sd391, 32'sd750,
32'sd744, 32'sd1235, 32'sd1172, 32'sd1149, 32'sd1827, 32'sd1622,
32'sd104, 32'sd995, 32'sd575, 32'sd1500, 32'sd847, 32'sd1411,
32'sd394, 32'sd1280, 32'sd383, 32'sd267, 32'sd1745, 32'sd240,
32'sd613, 32'sd1694, 32'sd1666, 32'sd1868, 32'sd1301, 32'sd1612,
32'sd1061, 32'sd161, 32'sd229, 32'sd655, 32'sd1335, 32'sd260,
32'sd506, 32'sd230, 32'sd1130, 32'sd1269, 32'sd1450, 32'sd1270,
32'sd894, 32'sd190, 32'sd1969, 32'sd1131, 32'sd998, 32'sd1904,
32'sd1992, 32'sd804, 32'sd1006, 32'sd1878, 32'sd104, 32'sd285,
32'sd378, 32'sd371, 32'sd1724, 32'sd1390, 32'sd1621, 32'sd1252,
32'sd1792, 32'sd1380, 32'sd1116, 32'sd438, 32'sd1868, 32'sd918,
32'sd1018, 32'sd205, 32'sd732, 32'sd1249, 32'sd1355, 32'sd1434,
32'sd220, 32'sd1629, 32'sd679, 32'sd764, 32'sd1748, 32'sd1192,
32'sd932, 32'sd1430, 32'sd394, 32'sd936, 32'sd1096, 32'sd511,
32'sd1741, 32'sd319, 32'sd1571, 32'sd945, 32'sd820, 32'sd272,
32'sd726, 32'sd1835, 32'sd1402, 32'sd596, 32'sd229, 32'sd1712,
32'sd529, 32'sd1061, 32'sd315, 32'sd1348, 32'sd1683, 32'sd1746,
32'sd1900, 32'sd1366, 32'sd1177, 32'sd1688, 32'sd1009, 32'sd1714,
32'sd710, 32'sd1526, 32'sd1219, 32'sd1545, 32'sd1534, 32'sd148,
32'sd1806, 32'sd1427, 32'sd1070, 32'sd1475, 32'sd1387, 32'sd629,
32'sd368, 32'sd1325, 32'sd511, 32'sd696, 32'sd1627, 32'sd706,
32'sd1305, 32'sd1747, 32'sd930, 32'sd1735, 32'sd1319, 32'sd1867,
32'sd188, 32'sd1259, 32'sd1180, 32'sd1348, 32'sd1949, 32'sd278,
32'sd614, 32'sd1539, 32'sd1387, 32'sd1575, 32'sd952, 32'sd822,
32'sd1793, 32'sd1569, 32'sd409, 32'sd275, 32'sd1719, 32'sd977,
32'sd864, 32'sd1325, 32'sd1200, 32'sd1539, 32'sd1640, 32'sd738,
32'sd294, 32'sd354, 32'sd1406, 32'sd1838, 32'sd762, 32'sd1639,
32'sd821, 32'sd343, 32'sd219, 32'sd1630, 32'sd108, 32'sd1664,
32'sd675, 32'sd983, 32'sd1304, 32'sd1350, 32'sd1066, 32'sd374,
32'sd1064, 32'sd1411, 32'sd339, 32'sd1232, 32'sd1215, 32'sd1952,
32'sd1987, 32'sd1339, 32'sd219, 32'sd1614, 32'sd1810, 32'sd1602,
32'sd1062, 32'sd1537, 32'sd868, 32'sd1644, 32'sd1789, 32'sd286,
32'sd837, 32'sd1795, 32'sd179, 32'sd191, 32'sd1601, 32'sd1578,
32'sd721, 32'sd1005, 32'sd1663, 32'sd1558, 32'sd1191, 32'sd753,
32'sd1906, 32'sd976, 32'sd1862, 32'sd1077, 32'sd1295, 32'sd1941,
32'sd640, 32'sd873, 32'sd1363, 32'sd1317, 32'sd1308, 32'sd1091,
32'sd482, 32'sd143, 32'sd261, 32'sd832, 32'sd1748, 32'sd223,
32'sd1935, 32'sd1198, 32'sd1171, 32'sd410, 32'sd321, 32'sd1172,
32'sd1029, 32'sd1095, 32'sd1285, 32'sd508, 32'sd704, 32'sd465,
32'sd1101, 32'sd1514, 32'sd1453, 32'sd1258, 32'sd1296, 32'sd397,
32'sd365, 32'sd862, 32'sd512, 32'sd329, 32'sd1390, 32'sd1625,
32'sd120, 32'sd778, 32'sd258, 32'sd1638, 32'sd177, 32'sd1721,
32'sd1503, 32'sd1943, 32'sd494, 32'sd948, 32'sd1877, 32'sd1356,
32'sd1880, 32'sd1912, 32'sd642, 32'sd1496, 32'sd409, 32'sd494,
32'sd1536, 32'sd1552, 32'sd933, 32'sd1317, 32'sd501, 32'sd190,
32'sd126, 32'sd1512, 32'sd468, 32'sd722, 32'sd277, 32'sd984,
32'sd306, 32'sd272, 32'sd1003, 32'sd1374, 32'sd1563, 32'sd319,
32'sd1542, 32'sd550, 32'sd1411, 32'sd1527, 32'sd480, 32'sd348,
32'sd1757, 32'sd1932, 32'sd1135, 32'sd1162, 32'sd844, 32'sd1081,
32'sd718, 32'sd1037, 32'sd714, 32'sd1282, 32'sd1690, 32'sd1848,
32'sd1162, 32'sd615, 32'sd1357, 32'sd362, 32'sd380, 32'sd343,
32'sd1002, 32'sd1772, 32'sd369, 32'sd781, 32'sd562, 32'sd422,
32'sd400, 32'sd851, 32'sd1759, 32'sd622, 32'sd724, 32'sd143,
32'sd204, 32'sd668, 32'sd1554, 32'sd1528, 32'sd1803, 32'sd1466,
32'sd1364, 32'sd162, 32'sd247, 32'sd1456, 32'sd1927, 32'sd1642,
32'sd1494, 32'sd563, 32'sd1672, 32'sd1959, 32'sd119, 32'sd1511,
32'sd855, 32'sd1423, 32'sd1342, 32'sd880, 32'sd1302, 32'sd386,
32'sd182, 32'sd1322, 32'sd238, 32'sd1226, 32'sd1919, 32'sd877,
32'sd463, 32'sd1384, 32'sd1868, 32'sd351, 32'sd165, 32'sd1626,
32'sd1229, 32'sd715, 32'sd450, 32'sd1748, 32'sd526, 32'sd845,
32'sd1987, 32'sd1692, 32'sd1490, 32'sd773, 32'sd1114, 32'sd1048,
32'sd1642, 32'sd376, 32'sd672, 32'sd1460, 32'sd1874, 32'sd1903,
32'sd650, 32'sd829, 32'sd748, 32'sd1159, 32'sd468, 32'sd907,
32'sd1933, 32'sd1158, 32'sd732, 32'sd609, 32'sd1267, 32'sd878,
32'sd1229, 32'sd419, 32'sd1329, 32'sd138, 32'sd1959, 32'sd1227,
32'sd1595, 32'sd1766, 32'sd1595, 32'sd1369, 32'sd1880, 32'sd263,
32'sd739, 32'sd769, 32'sd547, 32'sd295, 32'sd1251, 32'sd1213,
32'sd1338, 32'sd861, 32'sd915, 32'sd633, 32'sd1529, 32'sd1339,
32'sd982, 32'sd1886, 32'sd525, 32'sd937, 32'sd934, 32'sd1136,
32'sd570, 32'sd713, 32'sd554, 32'sd1865, 32'sd852, 32'sd1636,
32'sd1891, 32'sd1742, 32'sd1685, 32'sd1365, 32'sd1037, 32'sd1410,
32'sd1472, 32'sd518, 32'sd1871, 32'sd1455, 32'sd1273, 32'sd1872,
32'sd616, 32'sd924, 32'sd1065, 32'sd1679, 32'sd113, 32'sd502,
32'sd1416, 32'sd197, 32'sd1244, 32'sd821, 32'sd911, 32'sd1951,
32'sd128, 32'sd1323, 32'sd1899, 32'sd806, 32'sd746, 32'sd774,
32'sd1329, 32'sd1523, 32'sd255, 32'sd971, 32'sd663, 32'sd578,
32'sd1569, 32'sd1168, 32'sd769, 32'sd1119, 32'sd385, 32'sd112,
32'sd308, 32'sd1331, 32'sd1223, 32'sd1529, 32'sd1198, 32'sd845,
32'sd171, 32'sd841, 32'sd1665, 32'sd1004, 32'sd1989, 32'sd1282,
32'sd1788, 32'sd449, 32'sd175, 32'sd987, 32'sd1080, 32'sd263,
32'sd429, 32'sd1826, 32'sd156, 32'sd358, 32'sd978, 32'sd185,
32'sd295, 32'sd1386, 32'sd1747, 32'sd1590, 32'sd230, 32'sd374,
32'sd338, 32'sd476, 32'sd1611, 32'sd1635, 32'sd1461, 32'sd555,
32'sd458, 32'sd608, 32'sd722, 32'sd1393, 32'sd1534, 32'sd1254,
32'sd464, 32'sd1939, 32'sd1825, 32'sd1283, 32'sd1663, 32'sd1498,
32'sd312, 32'sd1679, 32'sd1701, 32'sd430, 32'sd1567, 32'sd655,
32'sd1884, 32'sd126, 32'sd292, 32'sd1498, 32'sd996, 32'sd503,
32'sd1403, 32'sd485, 32'sd211, 32'sd1001, 32'sd104, 32'sd745,
32'sd764, 32'sd986, 32'sd1497, 32'sd1853, 32'sd342, 32'sd1759,
32'sd1622, 32'sd587, 32'sd349, 32'sd1838, 32'sd1282, 32'sd1623,
32'sd307, 32'sd1294, 32'sd410, 32'sd627, 32'sd540, 32'sd428,
32'sd188, 32'sd829, 32'sd1472, 32'sd1738, 32'sd1145, 32'sd1055,
32'sd1903, 32'sd1553, 32'sd630, 32'sd438, 32'sd1118, 32'sd956,
32'sd296, 32'sd844, 32'sd1573, 32'sd1004, 32'sd1809, 32'sd1649,
32'sd1570, 32'sd1135, 32'sd1526, 32'sd184, 32'sd452, 32'sd119,
32'sd1232, 32'sd1142, 32'sd1892, 32'sd1310, 32'sd1580, 32'sd960,
32'sd1223, 32'sd1821, 32'sd637, 32'sd1690, 32'sd1245, 32'sd1302,
32'sd938, 32'sd469, 32'sd1159, 32'sd708, 32'sd190, 32'sd1799,
32'sd1612, 32'sd1855, 32'sd1467, 32'sd555, 32'sd1440, 32'sd841,
32'sd1679, 32'sd1420, 32'sd362, 32'sd904, 32'sd1908, 32'sd1635,
32'sd269, 32'sd636, 32'sd1398, 32'sd406, 32'sd1749, 32'sd1554,
32'sd1591, 32'sd806, 32'sd592, 32'sd1857, 32'sd626, 32'sd520,
32'sd1576, 32'sd1494, 32'sd1464, 32'sd603, 32'sd619, 32'sd1706,
32'sd1609, 32'sd1962, 32'sd735, 32'sd1398, 32'sd229, 32'sd601,
32'sd1525, 32'sd708, 32'sd998, 32'sd1513, 32'sd172, 32'sd689,
32'sd130, 32'sd1066, 32'sd933, 32'sd1129, 32'sd823, 32'sd146,
32'sd1273, 32'sd1770, 32'sd236, 32'sd130, 32'sd1781, 32'sd1660,
32'sd744, 32'sd256, 32'sd1462, 32'sd865, 32'sd212, 32'sd1979,
32'sd229, 32'sd1550, 32'sd734, 32'sd511, 32'sd1111, 32'sd444,
32'sd1398, 32'sd1532, 32'sd1608, 32'sd131, 32'sd258, 32'sd1693,
32'sd1708, 32'sd1071, 32'sd374, 32'sd539, 32'sd1472, 32'sd1499,
32'sd1975, 32'sd1685, 32'sd576, 32'sd1994, 32'sd1998, 32'sd1643,
32'sd625, 32'sd458, 32'sd741, 32'sd1217, 32'sd924, 32'sd592,
32'sd337, 32'sd1020, 32'sd643, 32'sd1484, 32'sd945, 32'sd1128,
32'sd733, 32'sd1590, 32'sd875, 32'sd1214, 32'sd210, 32'sd1425,
32'sd911, 32'sd1439, 32'sd368, 32'sd1197, 32'sd397, 32'sd1779,
32'sd552, 32'sd532, 32'sd362, 32'sd1320, 32'sd1787, 32'sd896,
32'sd364, 32'sd1528, 32'sd517, 32'sd1060, 32'sd698, 32'sd644,
32'sd1403, 32'sd1996, 32'sd217, 32'sd836, 32'sd1868, 32'sd1258,
32'sd385, 32'sd361, 32'sd1884, 32'sd182, 32'sd640, 32'sd1339,
32'sd1271, 32'sd307, 32'sd1741, 32'sd978, 32'sd384, 32'sd969,
32'sd154, 32'sd1213, 32'sd1012, 32'sd981, 32'sd315, 32'sd1972,
32'sd1399, 32'sd219, 32'sd1583, 32'sd1261, 32'sd900, 32'sd630,
32'sd1891, 32'sd388, 32'sd960, 32'sd641, 32'sd881, 32'sd423,
32'sd1101, 32'sd800, 32'sd1092, 32'sd1807, 32'sd1561, 32'sd1417,
32'sd468, 32'sd1142, 32'sd735, 32'sd555, 32'sd1026, 32'sd420,
32'sd662, 32'sd296, 32'sd336, 32'sd824, 32'sd1881, 32'sd1872,
32'sd316, 32'sd255, 32'sd386, 32'sd502, 32'sd854, 32'sd1731,
32'sd1727, 32'sd144, 32'sd1014, 32'sd856, 32'sd721, 32'sd1539,
32'sd832, 32'sd223, 32'sd160, 32'sd768, 32'sd505, 32'sd1970,
32'sd1021, 32'sd1228, 32'sd1293, 32'sd583, 32'sd838, 32'sd1218,
32'sd1164, 32'sd502, 32'sd872, 32'sd1599, 32'sd776, 32'sd1921,
32'sd1982, 32'sd1477, 32'sd1472, 32'sd1281, 32'sd123, 32'sd1247,
32'sd353, 32'sd1008, 32'sd618, 32'sd1074, 32'sd792, 32'sd1409,
32'sd1738, 32'sd387, 32'sd909, 32'sd106, 32'sd967, 32'sd1426,
32'sd820, 32'sd222, 32'sd1625, 32'sd1836, 32'sd1165, 32'sd229,
32'sd1071, 32'sd1267, 32'sd507, 32'sd572, 32'sd750, 32'sd125,
32'sd918, 32'sd168, 32'sd1400, 32'sd377, 32'sd1765, 32'sd1560,
32'sd1067, 32'sd1759, 32'sd428, 32'sd1516, 32'sd247, 32'sd1303,
32'sd1058, 32'sd1267, 32'sd556, 32'sd1547, 32'sd763, 32'sd1706,
32'sd991, 32'sd1846, 32'sd1479, 32'sd1130, 32'sd457, 32'sd394,
32'sd1760, 32'sd1506, 32'sd1227, 32'sd271, 32'sd1634, 32'sd1978,
32'sd1331, 32'sd1972, 32'sd334, 32'sd1078, 32'sd1440, 32'sd1028,
32'sd1113, 32'sd1472, 32'sd1749, 32'sd1131, 32'sd268, 32'sd1653,
32'sd834, 32'sd290, 32'sd339, 32'sd117, 32'sd1299, 32'sd1140,
32'sd817, 32'sd1008, 32'sd552, 32'sd1168, 32'sd680, 32'sd1044,
32'sd454, 32'sd994, 32'sd558, 32'sd1521, 32'sd683, 32'sd1960,
32'sd1049, 32'sd1917, 32'sd676, 32'sd252, 32'sd181, 32'sd233,
32'sd1731, 32'sd391, 32'sd206, 32'sd717, 32'sd243, 32'sd384,
32'sd1601, 32'sd1904, 32'sd1865, 32'sd161, 32'sd1598, 32'sd714,
32'sd924, 32'sd487, 32'sd1677, 32'sd1691, 32'sd1518, 32'sd1325,
32'sd383, 32'sd1539, 32'sd332, 32'sd1896, 32'sd1325, 32'sd762,
32'sd1560, 32'sd745, 32'sd435, 32'sd1341, 32'sd1838, 32'sd1014,
32'sd1999, 32'sd1405, 32'sd870, 32'sd631, 32'sd751, 32'sd669,
32'sd831, 32'sd1158, 32'sd1006, 32'sd1970, 32'sd1287, 32'sd1775,
32'sd877, 32'sd1548, 32'sd754, 32'sd1094, 32'sd1536, 32'sd1255,
32'sd812, 32'sd1233, 32'sd378, 32'sd435, 32'sd629, 32'sd809,
32'sd199, 32'sd1907, 32'sd765, 32'sd217, 32'sd337, 32'sd125,
32'sd291, 32'sd1076, 32'sd450, 32'sd1956, 32'sd563, 32'sd1507,
32'sd872, 32'sd399, 32'sd615, 32'sd1553, 32'sd1546, 32'sd1103,
32'sd160, 32'sd1560, 32'sd1963, 32'sd1882, 32'sd766, 32'sd1831,
32'sd1698, 32'sd1368, 32'sd941, 32'sd256, 32'sd927, 32'sd244,
32'sd849, 32'sd956, 32'sd1690, 32'sd1104, 32'sd1596, 32'sd425,
32'sd1259, 32'sd1256, 32'sd1652, 32'sd1337, 32'sd1166, 32'sd1550,
32'sd1034, 32'sd1369, 32'sd1505, 32'sd1931, 32'sd1943, 32'sd1879,
32'sd918, 32'sd1702, 32'sd1124, 32'sd1641, 32'sd1568, 32'sd1818,
32'sd828, 32'sd1294, 32'sd1498, 32'sd1019, 32'sd1409, 32'sd1290,
32'sd442, 32'sd1570, 32'sd1774, 32'sd204, 32'sd989, 32'sd1967,
32'sd1658, 32'sd292, 32'sd1155, 32'sd163, 32'sd1548, 32'sd1567,
32'sd838, 32'sd359, 32'sd418, 32'sd922, 32'sd1121, 32'sd292,
32'sd225, 32'sd1896, 32'sd1315, 32'sd1441, 32'sd1786, 32'sd1956,
32'sd197, 32'sd534, 32'sd438, 32'sd1826, 32'sd507, 32'sd282,
32'sd1066, 32'sd166, 32'sd1700, 32'sd213, 32'sd1115, 32'sd1339,
32'sd1250, 32'sd1851, 32'sd1143, 32'sd1194, 32'sd1729, 32'sd179,
32'sd232, 32'sd566, 32'sd539, 32'sd1189, 32'sd1310, 32'sd1858,
32'sd520, 32'sd1952, 32'sd363, 32'sd1707, 32'sd604, 32'sd1560,
32'sd1922, 32'sd1226, 32'sd209, 32'sd888, 32'sd658, 32'sd1409,
32'sd905, 32'sd344, 32'sd921, 32'sd154, 32'sd467, 32'sd1910,
32'sd1537, 32'sd1446, 32'sd799, 32'sd1343, 32'sd1240, 32'sd525,
32'sd788, 32'sd639, 32'sd896, 32'sd815, 32'sd1913, 32'sd1372,
32'sd1360, 32'sd253, 32'sd732, 32'sd1425, 32'sd319, 32'sd468,
32'sd654, 32'sd1590, 32'sd1988, 32'sd1844, 32'sd1774, 32'sd485,
32'sd1035, 32'sd1853, 32'sd298, 32'sd1407, 32'sd1242, 32'sd949,
32'sd1381, 32'sd1485, 32'sd823, 32'sd374, 32'sd271, 32'sd1747,
32'sd1741, 32'sd220, 32'sd1042, 32'sd1223, 32'sd1133, 32'sd377,
32'sd1775, 32'sd944, 32'sd185, 32'sd1492, 32'sd228, 32'sd1470,
32'sd527, 32'sd911, 32'sd1789, 32'sd550, 32'sd863, 32'sd1728,
32'sd648, 32'sd1565, 32'sd1184, 32'sd912, 32'sd461, 32'sd1016,
32'sd1751, 32'sd835, 32'sd1970, 32'sd1118, 32'sd251, 32'sd598,
32'sd1588, 32'sd1440, 32'sd301, 32'sd1901, 32'sd143, 32'sd566,
32'sd1751, 32'sd378, 32'sd323, 32'sd167, 32'sd522, 32'sd1303,
32'sd1126, 32'sd1999, 32'sd784, 32'sd1837, 32'sd1768, 32'sd1431,
32'sd1465, 32'sd492, 32'sd1873, 32'sd1732, 32'sd1885, 32'sd294,
32'sd890, 32'sd1263, 32'sd1917, 32'sd334, 32'sd1766, 32'sd1560,
32'sd579, 32'sd1999, 32'sd543, 32'sd101, 32'sd1342, 32'sd1687,
32'sd1350, 32'sd1378, 32'sd1683, 32'sd107, 32'sd113, 32'sd877,
32'sd419, 32'sd1723, 32'sd1629, 32'sd1760, 32'sd741, 32'sd137,
32'sd1011, 32'sd1446, 32'sd1700, 32'sd324, 32'sd1336, 32'sd1607,
32'sd173, 32'sd604, 32'sd1021, 32'sd939, 32'sd653, 32'sd224,
32'sd1097, 32'sd395, 32'sd691, 32'sd1811, 32'sd1712, 32'sd1228,
32'sd335, 32'sd2000, 32'sd1813, 32'sd1048, 32'sd1671, 32'sd1292,
32'sd1720, 32'sd1423, 32'sd1883, 32'sd1884, 32'sd1640, 32'sd1214,
32'sd1594, 32'sd675, 32'sd1016, 32'sd1292, 32'sd1852, 32'sd1590,
32'sd1822, 32'sd780, 32'sd174, 32'sd1245, 32'sd1459, 32'sd1381,
32'sd1758, 32'sd1816, 32'sd1552, 32'sd1007, 32'sd1657, 32'sd984,
32'sd1537, 32'sd1842, 32'sd482, 32'sd486, 32'sd1288, 32'sd760,
32'sd473, 32'sd1455, 32'sd1861, 32'sd1729, 32'sd1782, 32'sd850,
32'sd521, 32'sd1140, 32'sd551, 32'sd1526, 32'sd728, 32'sd188,
32'sd1962, 32'sd1461, 32'sd447, 32'sd575, 32'sd1060, 32'sd951,
32'sd905, 32'sd256, 32'sd1443, 32'sd300, 32'sd1949, 32'sd1156,
32'sd1003, 32'sd1519, 32'sd949, 32'sd421, 32'sd1088, 32'sd1223,
32'sd871, 32'sd1985, 32'sd1753, 32'sd881, 32'sd947, 32'sd1945,
32'sd202, 32'sd1529, 32'sd695, 32'sd953, 32'sd1814, 32'sd416,
32'sd1149, 32'sd1164, 32'sd1349, 32'sd451, 32'sd249, 32'sd732,
32'sd1988, 32'sd1861, 32'sd1926, 32'sd1986, 32'sd1427, 32'sd125,
32'sd954, 32'sd631, 32'sd178, 32'sd988, 32'sd276, 32'sd1443,
32'sd1998, 32'sd282, 32'sd1572, 32'sd103, 32'sd182, 32'sd1834,
32'sd1441, 32'sd1821, 32'sd873, 32'sd870, 32'sd1768, 32'sd225,
32'sd663, 32'sd1727, 32'sd1965, 32'sd1718, 32'sd870, 32'sd1377,
32'sd1880, 32'sd739, 32'sd1585, 32'sd1220, 32'sd1830, 32'sd924,
32'sd1462, 32'sd1825, 32'sd397, 32'sd1637, 32'sd1940, 32'sd941,
32'sd1681, 32'sd143, 32'sd1283, 32'sd392, 32'sd1216, 32'sd1729,
32'sd1994, 32'sd715, 32'sd541, 32'sd405, 32'sd1714, 32'sd1023,
32'sd881, 32'sd163, 32'sd925, 32'sd518, 32'sd1296, 32'sd1128,
32'sd1903, 32'sd235, 32'sd1522, 32'sd749, 32'sd315, 32'sd689,
32'sd1199, 32'sd1231, 32'sd1732, 32'sd1188, 32'sd1411, 32'sd1181,
32'sd1988, 32'sd1424, 32'sd125, 32'sd1115, 32'sd595, 32'sd1642,
32'sd1701, 32'sd1580, 32'sd1969, 32'sd938, 32'sd1637, 32'sd1376,
32'sd1976, 32'sd1908, 32'sd1117, 32'sd900, 32'sd305, 32'sd1151,
32'sd536, 32'sd1866, 32'sd1064, 32'sd1368, 32'sd990, 32'sd1523,
32'sd832, 32'sd1604, 32'sd1960, 32'sd1333, 32'sd493, 32'sd165,
32'sd776, 32'sd190, 32'sd1966, 32'sd1914, 32'sd1152, 32'sd561,
32'sd423, 32'sd1385, 32'sd1034, 32'sd1876, 32'sd1547, 32'sd1622,
32'sd838, 32'sd1179, 32'sd1147, 32'sd1175, 32'sd153, 32'sd207,
32'sd1359, 32'sd793, 32'sd352, 32'sd1440, 32'sd1804, 32'sd1565,
32'sd549, 32'sd507, 32'sd1537, 32'sd1012, 32'sd504, 32'sd1730,
32'sd1075, 32'sd639, 32'sd554, 32'sd1481, 32'sd718, 32'sd368,
32'sd965, 32'sd1865, 32'sd1434, 32'sd1785, 32'sd1702, 32'sd414,
32'sd126, 32'sd1457, 32'sd1258, 32'sd434, 32'sd1635, 32'sd400,
32'sd1686, 32'sd1495, 32'sd1276, 32'sd1863, 32'sd1644, 32'sd1771,
32'sd1271, 32'sd1242, 32'sd1754, 32'sd211, 32'sd1530, 32'sd1791,
32'sd929, 32'sd654, 32'sd578, 32'sd255, 32'sd1110, 32'sd1093,
32'sd678, 32'sd877, 32'sd1385, 32'sd1411, 32'sd222, 32'sd598,
32'sd466, 32'sd252, 32'sd241, 32'sd423, 32'sd234, 32'sd176,
32'sd1274, 32'sd769, 32'sd907, 32'sd787, 32'sd143, 32'sd282,
32'sd764, 32'sd739, 32'sd1998, 32'sd688, 32'sd1155, 32'sd600,
32'sd715, 32'sd1750, 32'sd118, 32'sd1254, 32'sd127, 32'sd297,
32'sd1030, 32'sd151, 32'sd1166, 32'sd783, 32'sd674, 32'sd695,
32'sd420, 32'sd945, 32'sd1810, 32'sd818, 32'sd171, 32'sd1328,
32'sd1757, 32'sd610, 32'sd1916, 32'sd1650, 32'sd1507, 32'sd1025,
32'sd1792, 32'sd763, 32'sd1553, 32'sd614, 32'sd1635, 32'sd1402,
32'sd1924, 32'sd561, 32'sd1911, 32'sd369, 32'sd1545, 32'sd951,
32'sd992, 32'sd1979, 32'sd621, 32'sd685, 32'sd1572, 32'sd1155,
32'sd1529, 32'sd1888, 32'sd527, 32'sd1328, 32'sd1179, 32'sd947,
32'sd262, 32'sd799, 32'sd1384, 32'sd1194, 32'sd1580, 32'sd199,
32'sd1400, 32'sd1113, 32'sd168, 32'sd516, 32'sd476, 32'sd1567,
32'sd1089, 32'sd788, 32'sd1529, 32'sd1189, 32'sd489, 32'sd327,
32'sd266, 32'sd1095, 32'sd914, 32'sd1289, 32'sd1100, 32'sd627,
32'sd250, 32'sd1661, 32'sd1306, 32'sd496, 32'sd835, 32'sd972,
32'sd396, 32'sd555, 32'sd449, 32'sd1254, 32'sd1241, 32'sd1556,
32'sd414, 32'sd1297, 32'sd1027, 32'sd961, 32'sd164, 32'sd352,
32'sd349, 32'sd1967, 32'sd757, 32'sd1488, 32'sd602, 32'sd584,
32'sd871, 32'sd1429, 32'sd557, 32'sd470, 32'sd366, 32'sd758,
32'sd407, 32'sd1760, 32'sd306, 32'sd1613, 32'sd1501, 32'sd477,
32'sd365, 32'sd641, 32'sd1706, 32'sd1822, 32'sd1648, 32'sd1108,
32'sd1208, 32'sd940, 32'sd1636, 32'sd913, 32'sd486, 32'sd940,
32'sd1941, 32'sd923, 32'sd516, 32'sd1581, 32'sd108, 32'sd1622,
32'sd922, 32'sd409, 32'sd372, 32'sd271, 32'sd1600, 32'sd1430,
32'sd672, 32'sd928, 32'sd227, 32'sd885, 32'sd418, 32'sd204,
32'sd1346, 32'sd1579, 32'sd788, 32'sd1051, 32'sd1118, 32'sd556,
32'sd1743, 32'sd1549, 32'sd1544, 32'sd785, 32'sd1967, 32'sd215,
32'sd568, 32'sd298, 32'sd747, 32'sd1128, 32'sd1025, 32'sd1872,
32'sd1818, 32'sd113, 32'sd1519, 32'sd587, 32'sd637, 32'sd671,
32'sd1106, 32'sd1657, 32'sd723, 32'sd476, 32'sd1541, 32'sd1307,
32'sd1503, 32'sd592, 32'sd1282, 32'sd1700, 32'sd1024, 32'sd262,
32'sd1166, 32'sd1285, 32'sd126, 32'sd1241, 32'sd1630, 32'sd347,
32'sd1628, 32'sd862, 32'sd1525, 32'sd1651, 32'sd555, 32'sd472,
32'sd1692, 32'sd146, 32'sd1469, 32'sd441, 32'sd173, 32'sd1312,
32'sd948, 32'sd191, 32'sd1863, 32'sd143, 32'sd628, 32'sd1889,
32'sd549, 32'sd1736, 32'sd1898, 32'sd1059, 32'sd719, 32'sd1703,
32'sd1275, 32'sd591, 32'sd302, 32'sd1351, 32'sd440, 32'sd197,
32'sd1172, 32'sd1991, 32'sd900, 32'sd1782, 32'sd1613, 32'sd1817,
32'sd273, 32'sd1835, 32'sd998, 32'sd1048, 32'sd315, 32'sd318,
32'sd1960, 32'sd1309, 32'sd1307, 32'sd1975, 32'sd1422, 32'sd1791,
32'sd999, 32'sd762, 32'sd1685, 32'sd1282, 32'sd680, 32'sd1078,
32'sd921, 32'sd395, 32'sd489, 32'sd1065, 32'sd1509, 32'sd460,
32'sd849, 32'sd594, 32'sd1217, 32'sd584, 32'sd1828, 32'sd1573,
32'sd305, 32'sd297, 32'sd1616, 32'sd1321, 32'sd1943, 32'sd364,
32'sd1407, 32'sd1403, 32'sd1285, 32'sd182, 32'sd1201, 32'sd342,
32'sd455, 32'sd756, 32'sd1157, 32'sd646, 32'sd1579, 32'sd1740,
32'sd639, 32'sd616, 32'sd1881, 32'sd836, 32'sd1563, 32'sd1805,
32'sd1440, 32'sd403, 32'sd1449, 32'sd848, 32'sd1785, 32'sd1878,
32'sd1394, 32'sd1451, 32'sd207, 32'sd1429, 32'sd1022, 32'sd776,
32'sd1321, 32'sd200, 32'sd1835, 32'sd662, 32'sd263, 32'sd1928,
32'sd151, 32'sd1286, 32'sd659, 32'sd1888, 32'sd552, 32'sd1091,
32'sd1160, 32'sd1014, 32'sd1685, 32'sd184, 32'sd210, 32'sd1823,
32'sd1367, 32'sd1995, 32'sd1365, 32'sd136, 32'sd1624, 32'sd927,
32'sd289, 32'sd1575, 32'sd694, 32'sd1350, 32'sd1171, 32'sd742,
32'sd361, 32'sd1599, 32'sd630, 32'sd621, 32'sd1501, 32'sd1577,
32'sd332, 32'sd1270, 32'sd166, 32'sd1805, 32'sd1518, 32'sd1218,
32'sd1865, 32'sd576, 32'sd1217, 32'sd1233, 32'sd958, 32'sd506,
32'sd1401, 32'sd1879, 32'sd125, 32'sd138, 32'sd366, 32'sd1081,
32'sd1936, 32'sd1117, 32'sd724, 32'sd857, 32'sd1798, 32'sd1550,
32'sd471, 32'sd1943, 32'sd1098, 32'sd760, 32'sd760, 32'sd1147,
32'sd1411, 32'sd1810, 32'sd351, 32'sd473, 32'sd564, 32'sd1412,
32'sd1800, 32'sd1997, 32'sd153, 32'sd1168, 32'sd971, 32'sd185,
32'sd1683, 32'sd1794, 32'sd1327, 32'sd579, 32'sd1512, 32'sd487,
32'sd991, 32'sd1496, 32'sd174, 32'sd337, 32'sd1141, 32'sd372,
32'sd1048, 32'sd496, 32'sd344, 32'sd1576, 32'sd1236, 32'sd260,
32'sd289, 32'sd672, 32'sd850, 32'sd1196, 32'sd908, 32'sd658,
32'sd351, 32'sd1572, 32'sd1439, 32'sd245, 32'sd1076, 32'sd1850,
32'sd1530, 32'sd597, 32'sd1448, 32'sd198, 32'sd255, 32'sd1773,
32'sd479, 32'sd1811, 32'sd1956, 32'sd1912, 32'sd767, 32'sd148,
32'sd1508, 32'sd382, 32'sd117, 32'sd1406, 32'sd1778, 32'sd1545,
32'sd800, 32'sd1905, 32'sd819, 32'sd667, 32'sd1733, 32'sd1086,
32'sd673, 32'sd980, 32'sd1216, 32'sd1084, 32'sd1875, 32'sd122,
32'sd1385, 32'sd1397, 32'sd631, 32'sd1385, 32'sd1603, 32'sd1577,
32'sd128, 32'sd526, 32'sd1314, 32'sd1540, 32'sd1579, 32'sd127,
32'sd1653, 32'sd1122, 32'sd1918, 32'sd737, 32'sd1070, 32'sd536,
32'sd305, 32'sd1924, 32'sd1091, 32'sd1472, 32'sd1722, 32'sd1119,
32'sd176, 32'sd893, 32'sd422, 32'sd1036, 32'sd1282, 32'sd160,
32'sd1367, 32'sd1686, 32'sd1708, 32'sd1957, 32'sd667, 32'sd1451,
32'sd1751, 32'sd158, 32'sd382, 32'sd1809, 32'sd1240, 32'sd897,
32'sd531, 32'sd1977, 32'sd951, 32'sd1893, 32'sd1951, 32'sd575,
32'sd1351, 32'sd1596, 32'sd1631, 32'sd860, 32'sd1070, 32'sd1501,
32'sd1550, 32'sd1174, 32'sd1690, 32'sd1765, 32'sd541, 32'sd1939,
32'sd258, 32'sd498, 32'sd1854, 32'sd1201, 32'sd1768, 32'sd1507,
32'sd1510, 32'sd610, 32'sd254, 32'sd1204, 32'sd1892, 32'sd715,
32'sd1407, 32'sd396, 32'sd867, 32'sd1431, 32'sd1342, 32'sd1796,
32'sd1368, 32'sd1696, 32'sd870, 32'sd705, 32'sd1897, 32'sd370,
32'sd554, 32'sd1632, 32'sd394, 32'sd562, 32'sd1166, 32'sd1745,
32'sd326, 32'sd543, 32'sd822, 32'sd1464, 32'sd294, 32'sd264,
32'sd1430, 32'sd1940, 32'sd275, 32'sd979, 32'sd876, 32'sd1596,
32'sd412, 32'sd1858, 32'sd218, 32'sd779, 32'sd626, 32'sd826,
32'sd1648, 32'sd1210, 32'sd1841, 32'sd1359, 32'sd1908, 32'sd346,
32'sd1065, 32'sd1960, 32'sd1218, 32'sd1452, 32'sd1049, 32'sd593,
32'sd343, 32'sd882, 32'sd507, 32'sd1872, 32'sd1661, 32'sd1952,
32'sd940, 32'sd687, 32'sd299, 32'sd654, 32'sd1973, 32'sd978,
32'sd1328, 32'sd136, 32'sd501, 32'sd1100, 32'sd1127, 32'sd1010,
32'sd466, 32'sd1179, 32'sd1030, 32'sd1554, 32'sd1362, 32'sd124,
32'sd1317, 32'sd1629, 32'sd1479, 32'sd1230, 32'sd1986, 32'sd1453,
32'sd785, 32'sd1078, 32'sd434, 32'sd637, 32'sd1533, 32'sd625,
32'sd849, 32'sd1019, 32'sd712, 32'sd328, 32'sd399, 32'sd517,
32'sd1952, 32'sd1890, 32'sd1312, 32'sd1944, 32'sd1798, 32'sd1085,
32'sd909, 32'sd378, 32'sd864, 32'sd1923, 32'sd1898, 32'sd249,
32'sd529, 32'sd861, 32'sd1239, 32'sd1155, 32'sd1153, 32'sd1357,
32'sd1995, 32'sd131, 32'sd296, 32'sd1011, 32'sd1215, 32'sd1273,
32'sd467, 32'sd905, 32'sd704, 32'sd789, 32'sd297, 32'sd1199,
32'sd1391, 32'sd784, 32'sd1428, 32'sd997, 32'sd519, 32'sd1803,
32'sd1806, 32'sd722, 32'sd661, 32'sd1420, 32'sd116, 32'sd1104,
32'sd485, 32'sd970, 32'sd1171, 32'sd748, 32'sd483, 32'sd538,
32'sd1467, 32'sd109, 32'sd957, 32'sd1500, 32'sd138, 32'sd990,
32'sd1852, 32'sd539, 32'sd699, 32'sd1253, 32'sd1998, 32'sd1194,
32'sd1024, 32'sd645, 32'sd1171, 32'sd1039, 32'sd1350, 32'sd1656,
32'sd468, 32'sd1327, 32'sd954, 32'sd1611, 32'sd260, 32'sd880,
32'sd377, 32'sd630, 32'sd190, 32'sd578, 32'sd1611, 32'sd981,
32'sd1729, 32'sd586, 32'sd1343, 32'sd1739, 32'sd233, 32'sd428,
32'sd915, 32'sd1576, 32'sd1213, 32'sd134, 32'sd1231, 32'sd774,
32'sd858, 32'sd1176, 32'sd1652, 32'sd383, 32'sd285, 32'sd748,
32'sd505, 32'sd1922, 32'sd1481, 32'sd1904, 32'sd1442, 32'sd1072,
32'sd1946, 32'sd1346, 32'sd474, 32'sd743, 32'sd422, 32'sd403,
32'sd859, 32'sd776, 32'sd1905, 32'sd1548, 32'sd1389, 32'sd899,
32'sd1823, 32'sd669, 32'sd1113, 32'sd504, 32'sd380, 32'sd1792,
32'sd262, 32'sd585, 32'sd1123, 32'sd668, 32'sd1475, 32'sd540,
32'sd1275, 32'sd1591, 32'sd1309, 32'sd549, 32'sd1198, 32'sd1797,
32'sd731, 32'sd1467, 32'sd754, 32'sd1686, 32'sd746, 32'sd929,
32'sd153, 32'sd267, 32'sd1251, 32'sd1991, 32'sd1978, 32'sd1992,
32'sd197, 32'sd164, 32'sd990, 32'sd370, 32'sd1935, 32'sd1097,
32'sd1465, 32'sd753, 32'sd1656, 32'sd386, 32'sd1350, 32'sd419,
32'sd1318, 32'sd144, 32'sd1796, 32'sd1362, 32'sd156, 32'sd1324,
32'sd368, 32'sd500, 32'sd162, 32'sd731, 32'sd1081, 32'sd1306,
32'sd337, 32'sd1072, 32'sd684, 32'sd1800, 32'sd559, 32'sd461,
32'sd202, 32'sd597, 32'sd1171, 32'sd626, 32'sd625, 32'sd1859,
32'sd1831, 32'sd460, 32'sd647, 32'sd371, 32'sd214, 32'sd1373,
32'sd1557, 32'sd1285, 32'sd1389, 32'sd333, 32'sd322, 32'sd1194,
32'sd1490, 32'sd883, 32'sd1328, 32'sd1059, 32'sd283, 32'sd962,
32'sd853, 32'sd108, 32'sd896, 32'sd1078, 32'sd907, 32'sd1433,
32'sd1406, 32'sd1899, 32'sd119, 32'sd407, 32'sd1975, 32'sd404,
32'sd1713, 32'sd336, 32'sd570, 32'sd1112, 32'sd1918, 32'sd227,
32'sd357, 32'sd287, 32'sd407, 32'sd992, 32'sd742, 32'sd1257,
32'sd1403, 32'sd1088, 32'sd552, 32'sd1911, 32'sd1994, 32'sd1446,
32'sd1347, 32'sd1879, 32'sd764, 32'sd1580, 32'sd890, 32'sd249,
32'sd453, 32'sd1845, 32'sd1107, 32'sd1150, 32'sd800, 32'sd1195,
32'sd1045, 32'sd1195, 32'sd1517, 32'sd1357, 32'sd420, 32'sd774,
32'sd280, 32'sd1291, 32'sd1274, 32'sd961, 32'sd476, 32'sd996,
32'sd909, 32'sd200, 32'sd940, 32'sd146, 32'sd151, 32'sd1417,
32'sd388, 32'sd1053, 32'sd313, 32'sd1033, 32'sd508, 32'sd679,
32'sd1317, 32'sd969, 32'sd970, 32'sd1632, 32'sd795, 32'sd1166,
32'sd762, 32'sd419, 32'sd912, 32'sd910, 32'sd1009, 32'sd134,
32'sd914, 32'sd1919, 32'sd2000, 32'sd1328, 32'sd977, 32'sd803,
32'sd785, 32'sd1440, 32'sd1804, 32'sd379, 32'sd753, 32'sd851,
32'sd1226, 32'sd1785, 32'sd1690, 32'sd1615, 32'sd1381, 32'sd1547,
32'sd818, 32'sd1803, 32'sd706, 32'sd1506, 32'sd1043, 32'sd1426,
32'sd1393, 32'sd1320, 32'sd1189, 32'sd1347, 32'sd538, 32'sd299,
32'sd1408, 32'sd201, 32'sd1749, 32'sd158, 32'sd309, 32'sd723,
32'sd708, 32'sd1043, 32'sd554, 32'sd1469, 32'sd1255, 32'sd1031,
32'sd579, 32'sd1761, 32'sd591, 32'sd1603, 32'sd1919, 32'sd1103,
32'sd1659, 32'sd223, 32'sd1843, 32'sd472, 32'sd1420, 32'sd1830,
32'sd461, 32'sd1348, 32'sd453, 32'sd1479, 32'sd488, 32'sd987,
32'sd1161, 32'sd962, 32'sd1523, 32'sd649, 32'sd1149, 32'sd1785,
32'sd504, 32'sd1455, 32'sd1292, 32'sd1137, 32'sd615, 32'sd1026,
32'sd845, 32'sd1351, 32'sd210, 32'sd1587, 32'sd756, 32'sd308,
32'sd183, 32'sd723, 32'sd880, 32'sd572, 32'sd1299, 32'sd1888,
32'sd1657, 32'sd449, 32'sd1475, 32'sd1874, 32'sd1351, 32'sd1008,
32'sd1751, 32'sd191, 32'sd1388, 32'sd1096, 32'sd669, 32'sd228,
32'sd1925, 32'sd1004, 32'sd678, 32'sd1352, 32'sd1993, 32'sd1549,
32'sd1249, 32'sd1435, 32'sd956, 32'sd1711, 32'sd1184, 32'sd993,
32'sd794, 32'sd681, 32'sd1154, 32'sd1735, 32'sd1107, 32'sd795,
32'sd1069, 32'sd1064, 32'sd1796, 32'sd727, 32'sd105, 32'sd1269,
32'sd1200, 32'sd1072, 32'sd136, 32'sd1718, 32'sd831, 32'sd1558,
32'sd1809, 32'sd1158, 32'sd1869, 32'sd440, 32'sd1496, 32'sd1889,
32'sd986, 32'sd1135, 32'sd1144, 32'sd699, 32'sd1540, 32'sd1352,
32'sd1381, 32'sd353, 32'sd1836, 32'sd1200, 32'sd895, 32'sd1387,
32'sd1296, 32'sd796, 32'sd1127, 32'sd1335, 32'sd1807, 32'sd792,
32'sd1124, 32'sd316, 32'sd884, 32'sd993, 32'sd1908, 32'sd993,
32'sd1536, 32'sd1832, 32'sd1206, 32'sd187, 32'sd772, 32'sd222,
32'sd1236, 32'sd1611, 32'sd1650, 32'sd536, 32'sd1136, 32'sd418,
32'sd1942, 32'sd1391, 32'sd1446, 32'sd674, 32'sd1864, 32'sd475,
32'sd1866, 32'sd957, 32'sd1082, 32'sd1051, 32'sd935, 32'sd1877,
32'sd1944, 32'sd438, 32'sd250, 32'sd1772, 32'sd217, 32'sd540,
32'sd1001, 32'sd1380, 32'sd1011, 32'sd1952, 32'sd1781, 32'sd1642,
32'sd1144, 32'sd1026, 32'sd1808, 32'sd1686, 32'sd1314, 32'sd1813,
32'sd1673, 32'sd1526, 32'sd1798, 32'sd648, 32'sd1847, 32'sd179,
32'sd253, 32'sd608, 32'sd1161, 32'sd1238, 32'sd1434, 32'sd1040,
32'sd1115, 32'sd847, 32'sd1596, 32'sd358, 32'sd371, 32'sd1211,
32'sd688, 32'sd123, 32'sd1197, 32'sd883, 32'sd827, 32'sd768,
32'sd101, 32'sd108, 32'sd355, 32'sd1967, 32'sd172, 32'sd912,
32'sd1525, 32'sd760, 32'sd899, 32'sd737, 32'sd822, 32'sd1900,
32'sd1080, 32'sd1477, 32'sd486, 32'sd1067, 32'sd1252, 32'sd1711,
32'sd1884, 32'sd550, 32'sd950, 32'sd913, 32'sd873, 32'sd271,
32'sd1945, 32'sd155, 32'sd990, 32'sd635, 32'sd589, 32'sd1270,
32'sd1130, 32'sd1542, 32'sd1829, 32'sd821, 32'sd1565, 32'sd1823,
32'sd683, 32'sd1348, 32'sd1882, 32'sd1493, 32'sd1681, 32'sd332,
32'sd1739, 32'sd911, 32'sd808, 32'sd823, 32'sd1482, 32'sd1153,
32'sd803, 32'sd1294, 32'sd1430, 32'sd1859, 32'sd1916, 32'sd1138,
32'sd1221, 32'sd1304, 32'sd1624, 32'sd345, 32'sd241, 32'sd1380,
32'sd549, 32'sd1799, 32'sd1113, 32'sd1188, 32'sd944, 32'sd1453,
32'sd1759, 32'sd1141, 32'sd149, 32'sd440, 32'sd1286, 32'sd1364,
32'sd1877, 32'sd1663, 32'sd1344, 32'sd883, 32'sd759, 32'sd469,
32'sd1656, 32'sd1881, 32'sd530, 32'sd481, 32'sd1497, 32'sd123,
32'sd1897, 32'sd1592, 32'sd653, 32'sd985, 32'sd671, 32'sd1152,
32'sd1026, 32'sd1935, 32'sd1206, 32'sd466, 32'sd524, 32'sd1533,
32'sd440, 32'sd1069, 32'sd1072, 32'sd1617, 32'sd1211, 32'sd1092,
32'sd950, 32'sd387, 32'sd450, 32'sd1753, 32'sd987, 32'sd1723,
32'sd1881, 32'sd691, 32'sd1837, 32'sd1074, 32'sd903, 32'sd986,
32'sd698, 32'sd578, 32'sd625, 32'sd223, 32'sd1580, 32'sd572,
32'sd637, 32'sd137, 32'sd799, 32'sd461, 32'sd749, 32'sd1594,
32'sd1973, 32'sd542, 32'sd856, 32'sd269, 32'sd260, 32'sd906,
32'sd490, 32'sd742, 32'sd154, 32'sd554, 32'sd628, 32'sd1488,
32'sd301, 32'sd1745, 32'sd104, 32'sd333, 32'sd293, 32'sd380,
32'sd1064, 32'sd1566, 32'sd1774, 32'sd639, 32'sd429, 32'sd1204,
32'sd1825, 32'sd521, 32'sd179, 32'sd1242, 32'sd602, 32'sd1900,
32'sd1069, 32'sd540, 32'sd608, 32'sd595, 32'sd686, 32'sd1270,
32'sd640, 32'sd1315, 32'sd168, 32'sd835, 32'sd424, 32'sd771,
32'sd918, 32'sd891, 32'sd244, 32'sd410, 32'sd1305, 32'sd736,
32'sd1322, 32'sd566, 32'sd696, 32'sd332, 32'sd778, 32'sd1251,
32'sd398, 32'sd181, 32'sd1043, 32'sd1736, 32'sd1229, 32'sd138,
32'sd694, 32'sd543, 32'sd1965, 32'sd1932, 32'sd946, 32'sd896,
32'sd1657, 32'sd961, 32'sd1605, 32'sd1573, 32'sd1330, 32'sd1877,
32'sd1420, 32'sd185, 32'sd105, 32'sd469, 32'sd512, 32'sd1448,
32'sd1124, 32'sd162, 32'sd272, 32'sd102, 32'sd1162, 32'sd1932,
32'sd871, 32'sd171, 32'sd1807, 32'sd1774, 32'sd510, 32'sd703,
32'sd1874, 32'sd1958, 32'sd1920, 32'sd1978, 32'sd429, 32'sd357,
32'sd1727, 32'sd1121, 32'sd1589, 32'sd665, 32'sd1954, 32'sd617,
32'sd1012, 32'sd749, 32'sd945, 32'sd1493, 32'sd587, 32'sd401,
32'sd122, 32'sd1462, 32'sd1601, 32'sd1837, 32'sd415, 32'sd832,
32'sd1787, 32'sd1829, 32'sd1363, 32'sd1648, 32'sd1584, 32'sd1756,
32'sd211, 32'sd396, 32'sd635, 32'sd446, 32'sd1300, 32'sd1650,
32'sd1926, 32'sd663, 32'sd1948, 32'sd1299, 32'sd285, 32'sd1257,
32'sd1386, 32'sd1481, 32'sd794, 32'sd1204, 32'sd1558, 32'sd777,
32'sd1157, 32'sd1419, 32'sd1586, 32'sd254, 32'sd169, 32'sd1865,
32'sd237, 32'sd1858, 32'sd824, 32'sd613, 32'sd373, 32'sd1749,
32'sd1582, 32'sd235, 32'sd1901, 32'sd1837, 32'sd1520, 32'sd342,
32'sd186, 32'sd556, 32'sd426, 32'sd244, 32'sd1019, 32'sd1921,
32'sd203, 32'sd1395, 32'sd147, 32'sd587, 32'sd1537, 32'sd1524,
32'sd887, 32'sd1187, 32'sd212, 32'sd601, 32'sd1400, 32'sd949,
32'sd1359, 32'sd1301, 32'sd1264, 32'sd610, 32'sd1266, 32'sd172,
32'sd150, 32'sd443, 32'sd1677, 32'sd587, 32'sd1887, 32'sd190,
32'sd702, 32'sd446, 32'sd782, 32'sd1456, 32'sd1330, 32'sd1691,
32'sd1357, 32'sd1135, 32'sd924, 32'sd725, 32'sd1530, 32'sd330,
32'sd922, 32'sd543, 32'sd118, 32'sd528, 32'sd1454, 32'sd625,
32'sd471, 32'sd993, 32'sd1024, 32'sd1779, 32'sd1543, 32'sd1605,
32'sd177, 32'sd1307, 32'sd1403, 32'sd826, 32'sd1224, 32'sd1990,
32'sd581, 32'sd103, 32'sd1668, 32'sd1790, 32'sd269, 32'sd1784,
32'sd1853, 32'sd947, 32'sd749, 32'sd994, 32'sd1795, 32'sd169,
32'sd600, 32'sd1887, 32'sd1912, 32'sd462, 32'sd749, 32'sd1057,
32'sd182, 32'sd1410, 32'sd232, 32'sd516, 32'sd578, 32'sd739,
32'sd1201, 32'sd801, 32'sd1203, 32'sd893, 32'sd1241, 32'sd1555,
32'sd1308, 32'sd376, 32'sd1792, 32'sd696, 32'sd1221, 32'sd1114,
32'sd1964, 32'sd154, 32'sd139, 32'sd186, 32'sd1484, 32'sd1555,
32'sd1530, 32'sd191, 32'sd1871, 32'sd1800, 32'sd343, 32'sd1096,
32'sd1714, 32'sd466, 32'sd1063, 32'sd1954, 32'sd1508, 32'sd1313,
32'sd1601, 32'sd1887, 32'sd511, 32'sd101, 32'sd156, 32'sd1493,
32'sd267, 32'sd908, 32'sd1108, 32'sd1489, 32'sd887, 32'sd1100,
32'sd1028, 32'sd459, 32'sd664, 32'sd1064, 32'sd1484, 32'sd1838,
32'sd771, 32'sd1478, 32'sd1259, 32'sd1457, 32'sd814, 32'sd1850,
32'sd1683, 32'sd1502, 32'sd533, 32'sd1256, 32'sd1073, 32'sd559,
32'sd1905, 32'sd1011, 32'sd1279, 32'sd849, 32'sd1055, 32'sd955,
32'sd1431, 32'sd296, 32'sd1646, 32'sd1823, 32'sd1884, 32'sd1480,
32'sd1332, 32'sd550, 32'sd1540, 32'sd983, 32'sd172, 32'sd1218,
32'sd1524, 32'sd1526, 32'sd1536, 32'sd1706, 32'sd1184, 32'sd1370,
32'sd500, 32'sd604, 32'sd1320, 32'sd326, 32'sd208, 32'sd788,
32'sd546, 32'sd782, 32'sd1523, 32'sd902, 32'sd278, 32'sd1867,
32'sd117, 32'sd436, 32'sd1561, 32'sd936, 32'sd119, 32'sd487,
32'sd1776, 32'sd1245, 32'sd960, 32'sd231, 32'sd1072, 32'sd1166,
32'sd989, 32'sd341, 32'sd1021, 32'sd1256, 32'sd1648, 32'sd1463,
32'sd1571, 32'sd168, 32'sd705, 32'sd1878, 32'sd1142, 32'sd1022,
32'sd1104, 32'sd544, 32'sd249, 32'sd555, 32'sd1612, 32'sd1294,
32'sd653, 32'sd454, 32'sd550, 32'sd220, 32'sd1573, 32'sd1624,
32'sd385, 32'sd486, 32'sd433, 32'sd1579, 32'sd1157, 32'sd215,
32'sd1947, 32'sd176, 32'sd302, 32'sd1703, 32'sd986, 32'sd293,
32'sd846, 32'sd1065, 32'sd1587, 32'sd1566, 32'sd268, 32'sd943,
32'sd1231, 32'sd1391, 32'sd528, 32'sd178, 32'sd1335, 32'sd198,
32'sd748, 32'sd754, 32'sd1800, 32'sd1465, 32'sd686, 32'sd611,
32'sd755, 32'sd1977, 32'sd1947, 32'sd347, 32'sd1079, 32'sd1601,
32'sd851, 32'sd1988, 32'sd1868, 32'sd992, 32'sd1670, 32'sd120,
32'sd1108, 32'sd1887, 32'sd1637, 32'sd969, 32'sd582, 32'sd383,
32'sd766, 32'sd475, 32'sd1441, 32'sd442, 32'sd226, 32'sd1990,
32'sd459, 32'sd1596, 32'sd1305, 32'sd112, 32'sd1975, 32'sd1945,
32'sd691, 32'sd1349, 32'sd231, 32'sd1073, 32'sd1641, 32'sd1382,
32'sd632, 32'sd270, 32'sd1150, 32'sd1364, 32'sd883, 32'sd1612,
32'sd1924, 32'sd1843, 32'sd509, 32'sd1824, 32'sd343, 32'sd966,
32'sd562, 32'sd128, 32'sd851, 32'sd1259, 32'sd1925, 32'sd1105,
32'sd1640, 32'sd1418, 32'sd1660, 32'sd579, 32'sd1818, 32'sd1298,
32'sd1095, 32'sd659, 32'sd1369, 32'sd1816, 32'sd307, 32'sd986,
32'sd1109, 32'sd1460, 32'sd571, 32'sd1906, 32'sd118, 32'sd962,
32'sd839, 32'sd204, 32'sd637, 32'sd846, 32'sd357, 32'sd1555,
32'sd1225, 32'sd1458, 32'sd456, 32'sd218, 32'sd1505, 32'sd1410,
32'sd1537, 32'sd1270, 32'sd1487, 32'sd1473, 32'sd1368, 32'sd1100,
32'sd219, 32'sd939, 32'sd1960, 32'sd349, 32'sd924, 32'sd938,
32'sd200, 32'sd1475, 32'sd367, 32'sd313, 32'sd279, 32'sd155,
32'sd963, 32'sd1804, 32'sd1940, 32'sd124, 32'sd955, 32'sd1723,
32'sd725, 32'sd1757, 32'sd1418, 32'sd391, 32'sd1517, 32'sd173,
32'sd1143, 32'sd594, 32'sd717, 32'sd185, 32'sd246, 32'sd1945,
32'sd1830, 32'sd1345, 32'sd1938, 32'sd1469, 32'sd892, 32'sd533,
32'sd1111, 32'sd821, 32'sd1481, 32'sd835, 32'sd233, 32'sd652,
32'sd1668, 32'sd407, 32'sd301, 32'sd1476, 32'sd563, 32'sd1326,
32'sd1689, 32'sd496, 32'sd1629, 32'sd813, 32'sd1369, 32'sd149,
32'sd1202, 32'sd762, 32'sd424, 32'sd563, 32'sd1760, 32'sd226,
32'sd583, 32'sd1506, 32'sd182, 32'sd390, 32'sd1773, 32'sd679,
32'sd1138, 32'sd1928, 32'sd1088, 32'sd104, 32'sd1386, 32'sd1948,
32'sd549, 32'sd564, 32'sd495, 32'sd125, 32'sd1424, 32'sd1150,
32'sd832, 32'sd276, 32'sd248, 32'sd1307, 32'sd239, 32'sd1681,
32'sd1513, 32'sd1947, 32'sd1087, 32'sd783, 32'sd169, 32'sd706,
32'sd1045, 32'sd473, 32'sd557, 32'sd1662, 32'sd636, 32'sd1693,
32'sd1937, 32'sd1272, 32'sd781, 32'sd538, 32'sd363, 32'sd1926,
32'sd1162, 32'sd949, 32'sd1493, 32'sd1357, 32'sd1821, 32'sd1338,
32'sd1447, 32'sd1151, 32'sd147, 32'sd1311, 32'sd934, 32'sd1498,
32'sd233, 32'sd1012, 32'sd686, 32'sd1055, 32'sd1277, 32'sd1386,
32'sd1466, 32'sd611, 32'sd775, 32'sd225, 32'sd875, 32'sd1766,
32'sd624, 32'sd1653, 32'sd764, 32'sd104, 32'sd896, 32'sd1960,
32'sd1000, 32'sd1460, 32'sd1724, 32'sd515, 32'sd589, 32'sd117,
32'sd1334, 32'sd981, 32'sd386, 32'sd1481, 32'sd345, 32'sd317,
32'sd1521, 32'sd1518, 32'sd1015, 32'sd880, 32'sd1878, 32'sd182,
32'sd1972, 32'sd356, 32'sd489, 32'sd1937, 32'sd302, 32'sd106,
32'sd811, 32'sd1540, 32'sd674, 32'sd556, 32'sd1761, 32'sd126,
32'sd494, 32'sd1363, 32'sd334, 32'sd1641, 32'sd1294, 32'sd656,
32'sd1903, 32'sd2000, 32'sd1238, 32'sd851, 32'sd1170, 32'sd745,
32'sd1060, 32'sd1472, 32'sd700, 32'sd186, 32'sd744, 32'sd1152,
32'sd963, 32'sd1581, 32'sd384, 32'sd689, 32'sd277, 32'sd679,
32'sd1067, 32'sd1929, 32'sd1313, 32'sd781, 32'sd526, 32'sd1151,
32'sd1916, 32'sd1619, 32'sd1323, 32'sd1464, 32'sd1892, 32'sd500,
32'sd520, 32'sd801, 32'sd1847, 32'sd1183, 32'sd327, 32'sd1131,
32'sd668, 32'sd868, 32'sd211, 32'sd1205, 32'sd1025, 32'sd369,
32'sd716, 32'sd1918, 32'sd1573, 32'sd1355, 32'sd291, 32'sd138,
32'sd1862, 32'sd1356, 32'sd1388, 32'sd170, 32'sd277, 32'sd707,
32'sd308, 32'sd1489, 32'sd1446, 32'sd1362, 32'sd1308, 32'sd140,
32'sd1784, 32'sd621, 32'sd1888, 32'sd1018, 32'sd1156, 32'sd787,
32'sd599, 32'sd580, 32'sd1219, 32'sd545, 32'sd302, 32'sd1716,
32'sd1024, 32'sd1875, 32'sd1058, 32'sd337, 32'sd1878, 32'sd142,
32'sd462, 32'sd267, 32'sd1851, 32'sd1970, 32'sd1993, 32'sd1015,
32'sd1143, 32'sd570, 32'sd1269, 32'sd861, 32'sd106, 32'sd1534,
32'sd114, 32'sd1309, 32'sd1543, 32'sd1505, 32'sd1118, 32'sd439,
32'sd1162, 32'sd761, 32'sd1251, 32'sd1648, 32'sd1540, 32'sd1443,
32'sd1899, 32'sd986, 32'sd1317, 32'sd1949, 32'sd1104, 32'sd1952,
32'sd683, 32'sd1193, 32'sd320, 32'sd1285, 32'sd331, 32'sd957,
32'sd673, 32'sd192, 32'sd2000, 32'sd1800, 32'sd1632, 32'sd1528,
32'sd365, 32'sd1887, 32'sd115, 32'sd309, 32'sd930, 32'sd1224,
32'sd1772, 32'sd310, 32'sd319, 32'sd1897, 32'sd1722, 32'sd1765,
32'sd1635, 32'sd1347, 32'sd959, 32'sd329, 32'sd1123, 32'sd607,
32'sd155, 32'sd1661, 32'sd441, 32'sd1516, 32'sd1036, 32'sd1714,
32'sd885, 32'sd1794, 32'sd1256, 32'sd1062, 32'sd1629, 32'sd265,
32'sd181, 32'sd574, 32'sd1243, 32'sd1122, 32'sd1546, 32'sd1050,
32'sd410, 32'sd480, 32'sd1661, 32'sd443, 32'sd728, 32'sd715,
32'sd298, 32'sd671, 32'sd442, 32'sd843, 32'sd659, 32'sd1523,
32'sd104, 32'sd1383, 32'sd517, 32'sd1579, 32'sd637, 32'sd1274,
32'sd764, 32'sd671, 32'sd1812, 32'sd409, 32'sd602, 32'sd887,
32'sd215, 32'sd756, 32'sd1490, 32'sd684, 32'sd409, 32'sd1846,
32'sd1905, 32'sd1736, 32'sd358, 32'sd617, 32'sd1463, 32'sd1979,
32'sd1976, 32'sd207, 32'sd1302, 32'sd1235, 32'sd1900, 32'sd740,
32'sd1006, 32'sd990, 32'sd1976, 32'sd1404, 32'sd829, 32'sd1326,
32'sd727, 32'sd191, 32'sd305, 32'sd1885, 32'sd482, 32'sd1006,
32'sd1676, 32'sd2000, 32'sd725, 32'sd737, 32'sd1467, 32'sd1773,
32'sd161, 32'sd912, 32'sd615, 32'sd1911, 32'sd1281, 32'sd523,
32'sd1460, 32'sd163, 32'sd730, 32'sd1924, 32'sd633, 32'sd1978,
32'sd384, 32'sd391, 32'sd1820, 32'sd1259, 32'sd569, 32'sd1986,
32'sd563, 32'sd190, 32'sd1618, 32'sd1174, 32'sd185, 32'sd1406,
32'sd941, 32'sd1073, 32'sd1125, 32'sd1696, 32'sd1771, 32'sd528,
32'sd289, 32'sd329, 32'sd774, 32'sd328, 32'sd1265, 32'sd831,
32'sd889, 32'sd1952, 32'sd501, 32'sd1630, 32'sd1808, 32'sd1049,
32'sd512, 32'sd283, 32'sd1683, 32'sd1076, 32'sd733, 32'sd850,
32'sd1695, 32'sd1858, 32'sd747, 32'sd1722, 32'sd554, 32'sd936,
32'sd1672, 32'sd187, 32'sd1762, 32'sd625, 32'sd140, 32'sd1181,
32'sd658, 32'sd1264, 32'sd336, 32'sd1772, 32'sd784, 32'sd1170,
32'sd1637, 32'sd1594, 32'sd1000, 32'sd1920, 32'sd298, 32'sd1231,
32'sd741, 32'sd972, 32'sd1677, 32'sd628, 32'sd926, 32'sd1429,
32'sd890, 32'sd1499, 32'sd442, 32'sd1724, 32'sd458, 32'sd549,
32'sd608, 32'sd1001, 32'sd1679, 32'sd688, 32'sd540, 32'sd1534,
32'sd218, 32'sd854, 32'sd599, 32'sd928, 32'sd1811, 32'sd928,
32'sd269, 32'sd170, 32'sd1442, 32'sd1350, 32'sd569, 32'sd924,
32'sd1788, 32'sd1152, 32'sd1314, 32'sd686, 32'sd912, 32'sd1962,
32'sd1475, 32'sd1207, 32'sd1718, 32'sd1453, 32'sd1843, 32'sd916,
32'sd859, 32'sd380, 32'sd357, 32'sd1362, 32'sd563, 32'sd1694,
32'sd1758, 32'sd514, 32'sd1099, 32'sd1841, 32'sd696, 32'sd628,
32'sd1909, 32'sd1802, 32'sd1564, 32'sd293, 32'sd492, 32'sd1291,
32'sd467, 32'sd1786, 32'sd293, 32'sd414, 32'sd849, 32'sd184,
32'sd1728, 32'sd966, 32'sd1313, 32'sd852, 32'sd1885, 32'sd1976,
32'sd944, 32'sd717, 32'sd1505, 32'sd189, 32'sd758, 32'sd1293,
32'sd883, 32'sd1225, 32'sd1067, 32'sd1554, 32'sd479, 32'sd497,
32'sd234, 32'sd1438, 32'sd908, 32'sd315, 32'sd1736, 32'sd1672,
32'sd523, 32'sd707, 32'sd1260, 32'sd1758, 32'sd1748, 32'sd1390,
32'sd516, 32'sd203, 32'sd703, 32'sd1832, 32'sd256, 32'sd1274,
32'sd924, 32'sd638, 32'sd1082, 32'sd555, 32'sd1710, 32'sd1411,
32'sd790, 32'sd1427, 32'sd399, 32'sd550, 32'sd1142, 32'sd1411,
32'sd972, 32'sd1356, 32'sd1926, 32'sd1730, 32'sd261, 32'sd334,
32'sd1630, 32'sd1332, 32'sd1350, 32'sd866, 32'sd243, 32'sd823,
32'sd1794, 32'sd469, 32'sd1424, 32'sd122, 32'sd1782, 32'sd1413,
32'sd615, 32'sd885, 32'sd597, 32'sd1953, 32'sd1030, 32'sd675,
32'sd1945, 32'sd1455, 32'sd634, 32'sd247, 32'sd1868, 32'sd1054,
32'sd1941, 32'sd802, 32'sd1173, 32'sd1965, 32'sd1217, 32'sd1489,
32'sd435, 32'sd216, 32'sd452, 32'sd1832, 32'sd501, 32'sd731,
32'sd1755, 32'sd307, 32'sd815, 32'sd223, 32'sd630, 32'sd1295,
32'sd1679, 32'sd809, 32'sd1783, 32'sd1403, 32'sd1072, 32'sd427,
32'sd1293, 32'sd1736, 32'sd384, 32'sd1283, 32'sd194, 32'sd1154,
32'sd1551, 32'sd397, 32'sd576, 32'sd1978, 32'sd118, 32'sd164,
32'sd668, 32'sd408, 32'sd1229, 32'sd1430, 32'sd166, 32'sd1191,
32'sd1036, 32'sd1374, 32'sd721, 32'sd1981, 32'sd775, 32'sd1463,
32'sd459, 32'sd861, 32'sd1135, 32'sd1080, 32'sd1400, 32'sd680,
32'sd720, 32'sd1582, 32'sd1990, 32'sd304, 32'sd1900, 32'sd840,
32'sd696, 32'sd653, 32'sd1301, 32'sd1861, 32'sd1752, 32'sd361,
32'sd1377, 32'sd1650, 32'sd891, 32'sd191, 32'sd956, 32'sd1676,
32'sd1334, 32'sd106, 32'sd381, 32'sd1582, 32'sd1428, 32'sd724,
32'sd606, 32'sd1065, 32'sd503, 32'sd1717, 32'sd365, 32'sd382,
32'sd1171, 32'sd411, 32'sd799, 32'sd1632, 32'sd929, 32'sd688,
32'sd1935, 32'sd1018, 32'sd876, 32'sd893, 32'sd725, 32'sd1962,
32'sd1775, 32'sd533, 32'sd1837, 32'sd1020, 32'sd1657, 32'sd536,
32'sd1356, 32'sd1576, 32'sd1852, 32'sd721, 32'sd738, 32'sd1364,
32'sd1952, 32'sd554, 32'sd269, 32'sd1433, 32'sd1258, 32'sd527,
32'sd647, 32'sd1383, 32'sd594, 32'sd869, 32'sd733, 32'sd919,
32'sd1334, 32'sd229, 32'sd146, 32'sd1689, 32'sd1030, 32'sd250,
32'sd793, 32'sd886, 32'sd972, 32'sd490, 32'sd1190, 32'sd341,
32'sd1232, 32'sd1845, 32'sd1080, 32'sd170, 32'sd582, 32'sd536,
32'sd1758, 32'sd775, 32'sd1575, 32'sd902, 32'sd164, 32'sd869,
32'sd908, 32'sd1404, 32'sd158, 32'sd351, 32'sd709, 32'sd504,
32'sd446, 32'sd1495, 32'sd1547, 32'sd1146, 32'sd560, 32'sd124,
32'sd1735, 32'sd1771, 32'sd1265, 32'sd318, 32'sd762, 32'sd1542,
32'sd1461, 32'sd1443, 32'sd1356, 32'sd1347, 32'sd1937, 32'sd1758,
32'sd460, 32'sd1036, 32'sd1897, 32'sd295, 32'sd1941, 32'sd1577,
32'sd948, 32'sd1816, 32'sd1485, 32'sd1561, 32'sd1058, 32'sd1764,
32'sd380, 32'sd1377, 32'sd554, 32'sd1858, 32'sd1154, 32'sd1429,
32'sd1170, 32'sd395, 32'sd1808, 32'sd844, 32'sd1315, 32'sd392,
32'sd1996, 32'sd1052, 32'sd1912, 32'sd1213, 32'sd1889, 32'sd1374,
32'sd1390, 32'sd1238, 32'sd1514, 32'sd1399, 32'sd1425, 32'sd418,
32'sd451, 32'sd1081, 32'sd255, 32'sd1945, 32'sd648, 32'sd1247,
32'sd1196, 32'sd411, 32'sd1711, 32'sd891, 32'sd1277, 32'sd806,
32'sd1361, 32'sd1583, 32'sd1075, 32'sd1453, 32'sd1878, 32'sd1242,
32'sd1065, 32'sd584, 32'sd496, 32'sd631, 32'sd449, 32'sd1535,
32'sd1826, 32'sd1991, 32'sd1831, 32'sd1318, 32'sd504, 32'sd1730,
32'sd679, 32'sd1376, 32'sd888, 32'sd994, 32'sd1400, 32'sd1660,
32'sd1003, 32'sd1925, 32'sd1779, 32'sd1618, 32'sd1946, 32'sd1029,
32'sd454, 32'sd1699, 32'sd1503, 32'sd742, 32'sd1061, 32'sd1461,
32'sd463, 32'sd1740, 32'sd1538, 32'sd1800, 32'sd1889, 32'sd609,
32'sd1007, 32'sd1611, 32'sd224, 32'sd594, 32'sd1164, 32'sd172,
32'sd1500, 32'sd1643, 32'sd1520, 32'sd1072, 32'sd866, 32'sd1522,
32'sd295, 32'sd1317, 32'sd1794, 32'sd144, 32'sd292, 32'sd1771,
32'sd1538, 32'sd590, 32'sd1845, 32'sd1902, 32'sd1338, 32'sd1808,
32'sd760, 32'sd573, 32'sd126, 32'sd1561, 32'sd1221, 32'sd1950,
32'sd1989, 32'sd1303, 32'sd622, 32'sd340, 32'sd1539, 32'sd1580,
32'sd898, 32'sd1667, 32'sd1025, 32'sd1756, 32'sd475, 32'sd1259,
32'sd1512, 32'sd1842, 32'sd1489, 32'sd318, 32'sd1905, 32'sd126,
32'sd1353, 32'sd449, 32'sd879, 32'sd1517, 32'sd1766, 32'sd329,
32'sd164, 32'sd1610, 32'sd273, 32'sd177, 32'sd1555, 32'sd1156,
32'sd1902, 32'sd372, 32'sd735, 32'sd1713, 32'sd857, 32'sd450,
32'sd1602, 32'sd177, 32'sd1134, 32'sd1795, 32'sd404, 32'sd1465,
32'sd329, 32'sd408, 32'sd1544, 32'sd564, 32'sd1724, 32'sd1743,
32'sd1674, 32'sd222, 32'sd1596, 32'sd471, 32'sd455, 32'sd623,
32'sd520, 32'sd1996, 32'sd1118, 32'sd850, 32'sd1161, 32'sd1429,
32'sd945, 32'sd546, 32'sd340, 32'sd1549, 32'sd1857, 32'sd433,
32'sd764, 32'sd1359, 32'sd149, 32'sd1207, 32'sd1015, 32'sd1342,
32'sd1493, 32'sd1261, 32'sd758, 32'sd539, 32'sd1727, 32'sd1663,
32'sd894, 32'sd400, 32'sd1385, 32'sd847, 32'sd943, 32'sd1132,
32'sd1875, 32'sd1441, 32'sd1491, 32'sd1337, 32'sd1075, 32'sd1615,
32'sd225, 32'sd805, 32'sd158, 32'sd508, 32'sd347, 32'sd1224,
32'sd271, 32'sd1243, 32'sd671, 32'sd1453, 32'sd690, 32'sd1725,
32'sd604, 32'sd459, 32'sd477, 32'sd384, 32'sd707, 32'sd1267,
32'sd1667, 32'sd1745, 32'sd1276, 32'sd144, 32'sd1516, 32'sd912,
32'sd1293, 32'sd1080, 32'sd585, 32'sd907, 32'sd894, 32'sd219,
32'sd758, 32'sd460, 32'sd1381, 32'sd1126, 32'sd167, 32'sd1435,
32'sd1085, 32'sd167, 32'sd223, 32'sd1879, 32'sd619, 32'sd1127,
32'sd643, 32'sd1174, 32'sd1225, 32'sd1040, 32'sd215, 32'sd1203,
32'sd1909, 32'sd1453, 32'sd875, 32'sd1083, 32'sd1885, 32'sd1674,
32'sd451, 32'sd925, 32'sd1853, 32'sd1149, 32'sd1476, 32'sd1398,
32'sd1349, 32'sd203, 32'sd1533, 32'sd1819, 32'sd1288, 32'sd357,
32'sd1218, 32'sd349, 32'sd866, 32'sd882, 32'sd1186, 32'sd1160,
32'sd1909, 32'sd257, 32'sd1115, 32'sd986, 32'sd1861, 32'sd1420,
32'sd1064, 32'sd445, 32'sd667, 32'sd407, 32'sd1687, 32'sd855,
32'sd1456, 32'sd1105, 32'sd1750, 32'sd1603, 32'sd1138, 32'sd244,
32'sd204, 32'sd1815, 32'sd1592, 32'sd306, 32'sd1766, 32'sd1939,
32'sd213, 32'sd1132, 32'sd124, 32'sd592, 32'sd362, 32'sd996,
32'sd828, 32'sd1637, 32'sd525, 32'sd1202, 32'sd1433, 32'sd1154,
32'sd1262, 32'sd1745, 32'sd1810, 32'sd630, 32'sd1742, 32'sd373,
32'sd1643, 32'sd992, 32'sd832, 32'sd991, 32'sd832, 32'sd1108,
32'sd1530, 32'sd935, 32'sd126, 32'sd1254, 32'sd276, 32'sd620,
32'sd490, 32'sd556, 32'sd1667, 32'sd308, 32'sd730, 32'sd995,
32'sd231, 32'sd1577, 32'sd725, 32'sd1890, 32'sd1592, 32'sd540,
32'sd1346, 32'sd620, 32'sd702, 32'sd1405, 32'sd517, 32'sd713,
32'sd1051, 32'sd1263, 32'sd1437, 32'sd250, 32'sd672, 32'sd365,
32'sd1492, 32'sd1411, 32'sd794, 32'sd370, 32'sd1219, 32'sd923,
32'sd1081, 32'sd1835, 32'sd202, 32'sd1884, 32'sd1894, 32'sd1238,
32'sd651, 32'sd1583, 32'sd1055, 32'sd204, 32'sd1730, 32'sd1329,
32'sd1579, 32'sd1462, 32'sd1160, 32'sd573, 32'sd1366, 32'sd612,
32'sd262, 32'sd511, 32'sd687, 32'sd953, 32'sd1508, 32'sd992,
32'sd1268, 32'sd1167, 32'sd955, 32'sd779, 32'sd1717, 32'sd1000,
32'sd1334, 32'sd578, 32'sd150, 32'sd571, 32'sd855, 32'sd587,
32'sd1063, 32'sd1983, 32'sd1330, 32'sd879, 32'sd1569, 32'sd1297,
32'sd1076, 32'sd673, 32'sd859, 32'sd427, 32'sd1119, 32'sd1082,
32'sd698, 32'sd775, 32'sd473, 32'sd1899, 32'sd1157, 32'sd612,
32'sd1828, 32'sd1275, 32'sd296, 32'sd217, 32'sd711, 32'sd843,
32'sd1189, 32'sd1815, 32'sd323, 32'sd1631, 32'sd468, 32'sd1188,
32'sd591, 32'sd479, 32'sd1638, 32'sd1774, 32'sd1122, 32'sd1568,
32'sd346, 32'sd1998, 32'sd1473, 32'sd1050, 32'sd1436, 32'sd1080,
32'sd140, 32'sd1756, 32'sd1426, 32'sd955, 32'sd113, 32'sd1078,
32'sd129, 32'sd565, 32'sd1632, 32'sd1814, 32'sd174, 32'sd708,
32'sd182, 32'sd943, 32'sd1690, 32'sd423, 32'sd1127, 32'sd1330,
32'sd1231, 32'sd949, 32'sd1514, 32'sd477, 32'sd852, 32'sd533,
32'sd1420, 32'sd429, 32'sd302, 32'sd1306, 32'sd1916, 32'sd1226,
32'sd1310, 32'sd443, 32'sd1949, 32'sd502, 32'sd633, 32'sd1976,
32'sd1119, 32'sd629, 32'sd874, 32'sd174, 32'sd582, 32'sd1233,
32'sd1334, 32'sd1875, 32'sd1738, 32'sd724, 32'sd1557, 32'sd1583,
32'sd668, 32'sd1568, 32'sd1186, 32'sd1682, 32'sd820, 32'sd881,
32'sd1461, 32'sd1111, 32'sd1865, 32'sd708, 32'sd340, 32'sd411,
32'sd1815, 32'sd454, 32'sd636, 32'sd224, 32'sd490, 32'sd130,
32'sd1200, 32'sd1124, 32'sd1496, 32'sd1229, 32'sd454, 32'sd966,
32'sd969, 32'sd937, 32'sd771, 32'sd1770, 32'sd923, 32'sd168,
32'sd613, 32'sd223, 32'sd696, 32'sd728, 32'sd1438, 32'sd567,
32'sd262, 32'sd930, 32'sd301, 32'sd1669, 32'sd1489, 32'sd877,
32'sd923, 32'sd698, 32'sd698, 32'sd692, 32'sd582, 32'sd1134,
32'sd1808, 32'sd1230, 32'sd174, 32'sd1219, 32'sd1141, 32'sd767,
32'sd1441, 32'sd745, 32'sd302, 32'sd1024, 32'sd295, 32'sd693,
32'sd448, 32'sd649, 32'sd691, 32'sd660, 32'sd362, 32'sd1665,
32'sd1462, 32'sd190, 32'sd817, 32'sd1948, 32'sd627, 32'sd431,
32'sd1145, 32'sd524, 32'sd1604, 32'sd1420, 32'sd438, 32'sd1736,
32'sd1230, 32'sd349, 32'sd649, 32'sd326, 32'sd638, 32'sd869,
32'sd1471, 32'sd1338, 32'sd1132, 32'sd306, 32'sd477, 32'sd1736,
32'sd1565, 32'sd1868, 32'sd253, 32'sd995, 32'sd178, 32'sd378,
32'sd109, 32'sd1112, 32'sd1300, 32'sd533, 32'sd1044, 32'sd470,
32'sd1308, 32'sd1574, 32'sd197, 32'sd1102, 32'sd168, 32'sd1939,
32'sd120, 32'sd752, 32'sd646, 32'sd1837, 32'sd583, 32'sd1248,
32'sd215, 32'sd951, 32'sd1904, 32'sd734, 32'sd1485, 32'sd1779,
32'sd1103, 32'sd628, 32'sd1010, 32'sd1373, 32'sd481, 32'sd242,
32'sd312, 32'sd413, 32'sd1472, 32'sd1989, 32'sd1788, 32'sd1252,
32'sd932, 32'sd469, 32'sd196, 32'sd1875, 32'sd449, 32'sd953,
32'sd731, 32'sd1926, 32'sd1737, 32'sd1598, 32'sd222, 32'sd1195,
32'sd796, 32'sd137, 32'sd1324, 32'sd523, 32'sd1674, 32'sd627,
32'sd836, 32'sd111, 32'sd1685, 32'sd1758, 32'sd692, 32'sd1326,
32'sd1761, 32'sd983, 32'sd1248, 32'sd1133, 32'sd1613, 32'sd1844,
32'sd710, 32'sd728, 32'sd1844, 32'sd1932, 32'sd1228, 32'sd1289,
32'sd447, 32'sd682, 32'sd1007, 32'sd1880, 32'sd847, 32'sd1866,
32'sd1371, 32'sd749, 32'sd1877, 32'sd1059, 32'sd1138, 32'sd1520,
32'sd1133, 32'sd1450, 32'sd147, 32'sd864, 32'sd1437, 32'sd405,
32'sd306, 32'sd1994, 32'sd238, 32'sd673, 32'sd1721, 32'sd824,
32'sd652, 32'sd205, 32'sd759, 32'sd1118, 32'sd407, 32'sd1917,
32'sd1607, 32'sd1898, 32'sd1611, 32'sd682, 32'sd1534, 32'sd1103,
32'sd862, 32'sd1214, 32'sd1028, 32'sd389, 32'sd753, 32'sd1809,
32'sd300, 32'sd1062, 32'sd1536, 32'sd1148, 32'sd1528, 32'sd202,
32'sd1590, 32'sd572, 32'sd1845, 32'sd1014, 32'sd516, 32'sd1440,
32'sd549, 32'sd1103, 32'sd399, 32'sd796, 32'sd624, 32'sd1132,
32'sd1876, 32'sd1802, 32'sd548, 32'sd1121, 32'sd1993, 32'sd930,
32'sd699, 32'sd120, 32'sd841, 32'sd890, 32'sd1057, 32'sd169,
32'sd929, 32'sd670, 32'sd1933, 32'sd446, 32'sd1334, 32'sd1499,
32'sd1447, 32'sd552, 32'sd1579, 32'sd1652, 32'sd1224, 32'sd101,
32'sd387, 32'sd698, 32'sd1857, 32'sd1605, 32'sd1297, 32'sd1355,
32'sd1021, 32'sd1697, 32'sd1539, 32'sd1850, 32'sd874, 32'sd177,
32'sd979, 32'sd1479, 32'sd484, 32'sd867, 32'sd745, 32'sd1261,
32'sd1711, 32'sd1657, 32'sd1952, 32'sd1994, 32'sd501, 32'sd253,
32'sd1030, 32'sd1319, 32'sd1557, 32'sd937, 32'sd1533, 32'sd1880,
32'sd937, 32'sd1015, 32'sd1880, 32'sd1133, 32'sd564, 32'sd410,
32'sd1321, 32'sd578, 32'sd1695, 32'sd1472, 32'sd786, 32'sd634,
32'sd1737, 32'sd1906, 32'sd376, 32'sd593, 32'sd1608, 32'sd1446,
32'sd980, 32'sd1061, 32'sd145, 32'sd1150, 32'sd1106, 32'sd1988,
32'sd1803, 32'sd671, 32'sd470, 32'sd906, 32'sd1267, 32'sd526,
32'sd768, 32'sd291, 32'sd830, 32'sd1061, 32'sd1964, 32'sd1707,
32'sd1395, 32'sd256, 32'sd1348, 32'sd1506, 32'sd1177, 32'sd301,
32'sd1874, 32'sd1237, 32'sd1483, 32'sd1544, 32'sd246, 32'sd1585,
32'sd1260, 32'sd1711, 32'sd411, 32'sd1118, 32'sd1878, 32'sd838,
32'sd212, 32'sd1325, 32'sd1295, 32'sd229, 32'sd251, 32'sd1499,
32'sd1597, 32'sd769, 32'sd1143, 32'sd652, 32'sd1519, 32'sd1747,
32'sd1647, 32'sd201, 32'sd530, 32'sd1109, 32'sd1599, 32'sd1388,
32'sd864, 32'sd727, 32'sd1428, 32'sd573, 32'sd160, 32'sd824,
32'sd722, 32'sd431, 32'sd823, 32'sd626, 32'sd565, 32'sd1898,
32'sd951, 32'sd1493, 32'sd1280, 32'sd1178, 32'sd271, 32'sd1751,
32'sd1568, 32'sd1565, 32'sd1405, 32'sd728, 32'sd893, 32'sd1466,
32'sd933, 32'sd592, 32'sd242, 32'sd1124, 32'sd1777, 32'sd575,
32'sd1891, 32'sd1796, 32'sd659, 32'sd1531, 32'sd1046, 32'sd161,
32'sd1368, 32'sd374, 32'sd1576, 32'sd1012, 32'sd1109, 32'sd1370,
32'sd1599, 32'sd1449, 32'sd1143, 32'sd1831, 32'sd1118, 32'sd1491,
32'sd1892, 32'sd1684, 32'sd1946, 32'sd989, 32'sd818, 32'sd1132,
32'sd435, 32'sd1649, 32'sd1984, 32'sd581, 32'sd690, 32'sd1009,
32'sd1871, 32'sd1889, 32'sd957, 32'sd1541, 32'sd701, 32'sd409,
32'sd1675, 32'sd1000, 32'sd386, 32'sd1278, 32'sd866, 32'sd1670,
32'sd279, 32'sd547, 32'sd182, 32'sd434, 32'sd1713, 32'sd1196,
32'sd220, 32'sd254, 32'sd1846, 32'sd151, 32'sd1104, 32'sd1562,
32'sd1628, 32'sd611, 32'sd385, 32'sd860, 32'sd1475, 32'sd523,
32'sd1534, 32'sd1855, 32'sd1338, 32'sd223, 32'sd1536, 32'sd1223,
32'sd1230, 32'sd1434, 32'sd1948, 32'sd1449, 32'sd204, 32'sd450,
32'sd1654, 32'sd1522, 32'sd1246, 32'sd818, 32'sd651, 32'sd1477,
32'sd1981, 32'sd1074, 32'sd1615, 32'sd863, 32'sd629, 32'sd392,
32'sd747, 32'sd865, 32'sd1046, 32'sd1390, 32'sd754, 32'sd872,
32'sd552, 32'sd931, 32'sd1774, 32'sd1798, 32'sd762, 32'sd756,
32'sd1970, 32'sd1333, 32'sd993, 32'sd1010, 32'sd293, 32'sd839,
32'sd994, 32'sd117, 32'sd664, 32'sd545, 32'sd1816, 32'sd1680,
32'sd480, 32'sd1438, 32'sd1979, 32'sd1105, 32'sd540, 32'sd1412,
32'sd572, 32'sd352, 32'sd473, 32'sd1148, 32'sd1947, 32'sd1527,
32'sd168, 32'sd1657, 32'sd860, 32'sd1095, 32'sd998, 32'sd1552,
32'sd1543, 32'sd457, 32'sd1131, 32'sd1605, 32'sd910, 32'sd101,
32'sd585, 32'sd1658, 32'sd274, 32'sd1097, 32'sd1558, 32'sd371,
32'sd865, 32'sd456, 32'sd743, 32'sd1902, 32'sd1392, 32'sd1840,
32'sd1166, 32'sd1964, 32'sd980, 32'sd511, 32'sd820, 32'sd852,
32'sd755, 32'sd224, 32'sd1377, 32'sd1374, 32'sd1348, 32'sd196,
32'sd1918, 32'sd864, 32'sd1391, 32'sd329, 32'sd870, 32'sd636,
32'sd1308, 32'sd1532, 32'sd1603, 32'sd315, 32'sd817, 32'sd330,
32'sd1771, 32'sd1239, 32'sd1235, 32'sd1238, 32'sd1928, 32'sd1161,
32'sd909, 32'sd1365, 32'sd393, 32'sd1446, 32'sd1548, 32'sd1595,
32'sd394, 32'sd1263, 32'sd1940, 32'sd723, 32'sd1746, 32'sd1338,
32'sd831, 32'sd1164, 32'sd246, 32'sd731, 32'sd1425, 32'sd1182,
32'sd1780, 32'sd1002, 32'sd1590, 32'sd856, 32'sd894, 32'sd1451,
32'sd1123, 32'sd1844, 32'sd906, 32'sd348, 32'sd903, 32'sd641,
32'sd1506, 32'sd937, 32'sd1003, 32'sd1722, 32'sd1026, 32'sd401,
32'sd637, 32'sd1698, 32'sd420, 32'sd329, 32'sd118, 32'sd1410,
32'sd157, 32'sd598, 32'sd1472, 32'sd670, 32'sd438, 32'sd1172,
32'sd896, 32'sd565, 32'sd134, 32'sd761, 32'sd1244, 32'sd157,
32'sd1849, 32'sd708, 32'sd1104, 32'sd1992, 32'sd1666, 32'sd194,
32'sd835, 32'sd1372, 32'sd1588, 32'sd1742, 32'sd1511, 32'sd1408,
32'sd434, 32'sd712, 32'sd1928, 32'sd1674, 32'sd251, 32'sd1564,
32'sd105, 32'sd1807, 32'sd1572, 32'sd925, 32'sd654, 32'sd1531,
32'sd427, 32'sd1406, 32'sd1799, 32'sd1956, 32'sd625, 32'sd950,
32'sd277, 32'sd1729, 32'sd1397, 32'sd679, 32'sd1212, 32'sd289,
32'sd871, 32'sd1249, 32'sd1308, 32'sd730, 32'sd1970, 32'sd947,
32'sd251, 32'sd356, 32'sd279, 32'sd531, 32'sd936, 32'sd664,
32'sd1192, 32'sd1695, 32'sd984, 32'sd225, 32'sd1399, 32'sd1918,
32'sd921, 32'sd1246, 32'sd1347, 32'sd970, 32'sd1626, 32'sd1420,
32'sd311, 32'sd1126, 32'sd1830, 32'sd1158, 32'sd429, 32'sd222,
32'sd900, 32'sd1989, 32'sd1978, 32'sd692, 32'sd612, 32'sd1878,
32'sd1314, 32'sd444, 32'sd979, 32'sd1951, 32'sd290, 32'sd1429,
32'sd1274, 32'sd1179, 32'sd1809, 32'sd1942, 32'sd523, 32'sd1558,
32'sd916, 32'sd355, 32'sd146, 32'sd407, 32'sd1285, 32'sd1669,
32'sd1836, 32'sd1919, 32'sd1410, 32'sd1140, 32'sd1333, 32'sd1201,
32'sd1776, 32'sd230, 32'sd1442, 32'sd1039, 32'sd282, 32'sd1218,
32'sd1868, 32'sd1710, 32'sd510, 32'sd946, 32'sd1715, 32'sd1299,
32'sd759, 32'sd1101, 32'sd1371, 32'sd648, 32'sd1520, 32'sd1214,
32'sd720, 32'sd997, 32'sd1762, 32'sd1843, 32'sd1699, 32'sd1431,
32'sd357, 32'sd305, 32'sd1889, 32'sd694, 32'sd1463, 32'sd1676,
32'sd1535, 32'sd677, 32'sd595, 32'sd776, 32'sd1866, 32'sd149,
32'sd1247, 32'sd627, 32'sd1269, 32'sd1845, 32'sd1176, 32'sd1611,
32'sd556, 32'sd810, 32'sd240, 32'sd1606, 32'sd267, 32'sd1299,
32'sd1584, 32'sd1999, 32'sd1386, 32'sd1804, 32'sd832, 32'sd534,
32'sd1519, 32'sd257, 32'sd571, 32'sd1583, 32'sd291, 32'sd1527,
32'sd1186, 32'sd1730, 32'sd1542, 32'sd1884, 32'sd1954, 32'sd144,
32'sd1130, 32'sd727, 32'sd758, 32'sd1083, 32'sd568, 32'sd482,
32'sd1454, 32'sd381, 32'sd100, 32'sd831, 32'sd212, 32'sd817,
32'sd1062, 32'sd1244, 32'sd1530, 32'sd1012, 32'sd984, 32'sd1079,
32'sd331, 32'sd946, 32'sd1392, 32'sd908, 32'sd851, 32'sd1820,
32'sd1990, 32'sd1204, 32'sd626, 32'sd882, 32'sd440, 32'sd1121,
32'sd800, 32'sd152, 32'sd1799, 32'sd187, 32'sd937, 32'sd684,
32'sd462, 32'sd1132, 32'sd1653, 32'sd1639, 32'sd1757, 32'sd662,
32'sd319, 32'sd981, 32'sd1249, 32'sd430, 32'sd868, 32'sd850,
32'sd701, 32'sd980, 32'sd1111, 32'sd488, 32'sd1910, 32'sd722,
32'sd1095, 32'sd1945, 32'sd137, 32'sd417, 32'sd493, 32'sd520,
32'sd1403, 32'sd655, 32'sd1036, 32'sd1616, 32'sd1953, 32'sd1105,
32'sd1109, 32'sd1835, 32'sd1088, 32'sd627, 32'sd1234, 32'sd284,
32'sd1725, 32'sd1438, 32'sd677, 32'sd708, 32'sd278, 32'sd1414,
32'sd596, 32'sd468, 32'sd1585, 32'sd1996, 32'sd141, 32'sd1282,
32'sd1317, 32'sd461, 32'sd1433, 32'sd1694, 32'sd961, 32'sd923,
32'sd1936, 32'sd680, 32'sd651, 32'sd340, 32'sd262, 32'sd345,
32'sd1974, 32'sd858, 32'sd584, 32'sd1526, 32'sd1024, 32'sd607,
32'sd1613, 32'sd1512, 32'sd549, 32'sd626, 32'sd495, 32'sd1868,
32'sd535, 32'sd1569, 32'sd254, 32'sd1018, 32'sd975, 32'sd1469,
32'sd463, 32'sd1922, 32'sd1519, 32'sd818, 32'sd547, 32'sd940,
32'sd1425, 32'sd1382, 32'sd544, 32'sd1047, 32'sd1249, 32'sd794,
32'sd170, 32'sd1872, 32'sd386, 32'sd1986, 32'sd807, 32'sd838,
32'sd171, 32'sd638, 32'sd1769, 32'sd203, 32'sd653, 32'sd397,
32'sd1255, 32'sd1283, 32'sd148, 32'sd703, 32'sd1368, 32'sd272,
32'sd268, 32'sd979, 32'sd1355, 32'sd1654, 32'sd1737, 32'sd951,
32'sd1175, 32'sd1991, 32'sd1828, 32'sd1026, 32'sd1687, 32'sd1436,
32'sd781, 32'sd494, 32'sd1020, 32'sd144, 32'sd1733, 32'sd1232,
32'sd1122, 32'sd1715, 32'sd457, 32'sd1354, 32'sd200, 32'sd100,
32'sd630, 32'sd527, 32'sd1347, 32'sd1836, 32'sd634, 32'sd1850,
32'sd1072, 32'sd1014, 32'sd1021, 32'sd1328, 32'sd463, 32'sd1312,
32'sd466, 32'sd551, 32'sd1966, 32'sd985, 32'sd1895, 32'sd1033,
32'sd221, 32'sd1025, 32'sd952, 32'sd904, 32'sd410, 32'sd1438,
32'sd2000, 32'sd1710, 32'sd555, 32'sd1338, 32'sd275, 32'sd1170,
32'sd1112, 32'sd951, 32'sd1021, 32'sd370, 32'sd892, 32'sd1585,
32'sd752, 32'sd683, 32'sd217, 32'sd742, 32'sd376, 32'sd1442,
32'sd1698, 32'sd1158, 32'sd906, 32'sd461, 32'sd1273, 32'sd665,
32'sd1485, 32'sd1797, 32'sd1368, 32'sd148, 32'sd1891, 32'sd299,
32'sd542, 32'sd390, 32'sd1186, 32'sd1335, 32'sd1401, 32'sd1377,
32'sd1200, 32'sd1981, 32'sd189, 32'sd107, 32'sd268, 32'sd1423,
32'sd102, 32'sd1141, 32'sd1942, 32'sd1029, 32'sd1699, 32'sd200,
32'sd1976, 32'sd939, 32'sd1547, 32'sd1807, 32'sd1488, 32'sd475,
32'sd1239, 32'sd287, 32'sd1435, 32'sd1503, 32'sd902, 32'sd825,
32'sd710, 32'sd1410, 32'sd1658, 32'sd189, 32'sd240, 32'sd759,
32'sd123, 32'sd1362, 32'sd576, 32'sd1153, 32'sd870, 32'sd1942,
32'sd1438, 32'sd568, 32'sd121, 32'sd781, 32'sd1823, 32'sd1376,
32'sd881, 32'sd1147, 32'sd362, 32'sd491, 32'sd996, 32'sd1080,
32'sd1214, 32'sd653, 32'sd1763, 32'sd916, 32'sd895, 32'sd1328,
32'sd1817, 32'sd219, 32'sd1675, 32'sd209, 32'sd1607, 32'sd1997,
32'sd363, 32'sd928, 32'sd140, 32'sd1369, 32'sd1934, 32'sd938,
32'sd280, 32'sd117, 32'sd1410, 32'sd747, 32'sd1683, 32'sd1229,
32'sd476, 32'sd1645, 32'sd1833, 32'sd1849, 32'sd1902, 32'sd1296,
32'sd860, 32'sd1795, 32'sd767, 32'sd206, 32'sd1216, 32'sd164,
32'sd1525, 32'sd1332, 32'sd1789, 32'sd720, 32'sd1517, 32'sd1884,
32'sd1199, 32'sd368, 32'sd604, 32'sd873, 32'sd1285, 32'sd672,
32'sd1342, 32'sd1340, 32'sd133, 32'sd1605, 32'sd227, 32'sd297,
32'sd515, 32'sd1998, 32'sd1987, 32'sd395, 32'sd1733, 32'sd994,
32'sd1974, 32'sd1392, 32'sd587, 32'sd261, 32'sd100, 32'sd665,
32'sd266, 32'sd475, 32'sd1313, 32'sd1038, 32'sd1162, 32'sd1306,
32'sd221, 32'sd506, 32'sd1619, 32'sd1552, 32'sd1185, 32'sd633,
32'sd1223, 32'sd1090, 32'sd720, 32'sd1093, 32'sd1191, 32'sd722,
32'sd894, 32'sd1130, 32'sd1191, 32'sd915, 32'sd1674, 32'sd274,
32'sd282, 32'sd843, 32'sd1009, 32'sd424, 32'sd1623, 32'sd1943,
32'sd933, 32'sd1431, 32'sd936, 32'sd800, 32'sd218, 32'sd1593,
32'sd1474, 32'sd1907, 32'sd626, 32'sd979, 32'sd210, 32'sd1515,
32'sd1986, 32'sd1941, 32'sd497, 32'sd949, 32'sd225, 32'sd1405,
32'sd1987, 32'sd156, 32'sd507, 32'sd1689, 32'sd1719, 32'sd655,
32'sd571, 32'sd1296, 32'sd1244, 32'sd610, 32'sd274, 32'sd674,
32'sd1732, 32'sd1752, 32'sd500, 32'sd1737, 32'sd1646, 32'sd609,
32'sd1050, 32'sd1077, 32'sd963, 32'sd471, 32'sd1740, 32'sd1176,
32'sd1245, 32'sd719, 32'sd1640, 32'sd1545, 32'sd698, 32'sd1000,
32'sd989, 32'sd1145, 32'sd1506, 32'sd124, 32'sd1442, 32'sd1983,
32'sd1666, 32'sd288, 32'sd1676, 32'sd1639, 32'sd660, 32'sd1042,
32'sd121, 32'sd896, 32'sd1248, 32'sd738, 32'sd1151, 32'sd1493,
32'sd1641, 32'sd1473, 32'sd1084, 32'sd1965, 32'sd1448, 32'sd819,
32'sd1818, 32'sd1154, 32'sd1633, 32'sd147, 32'sd222, 32'sd1252,
32'sd207, 32'sd1101, 32'sd1764, 32'sd1797, 32'sd1394, 32'sd1020,
32'sd1135, 32'sd1781, 32'sd956, 32'sd1857, 32'sd1285, 32'sd736,
32'sd874, 32'sd634, 32'sd678, 32'sd977, 32'sd1986, 32'sd1473,
32'sd276, 32'sd633, 32'sd778, 32'sd577, 32'sd1469, 32'sd1795,
32'sd1323, 32'sd587, 32'sd1201, 32'sd1328, 32'sd597, 32'sd947,
32'sd1555, 32'sd521, 32'sd355, 32'sd1243, 32'sd1361, 32'sd829,
32'sd1813, 32'sd266, 32'sd885, 32'sd1507, 32'sd1180, 32'sd1792,
32'sd1037, 32'sd1109, 32'sd1548, 32'sd1769, 32'sd1451, 32'sd464,
32'sd1311, 32'sd763, 32'sd788, 32'sd768, 32'sd368, 32'sd1892,
32'sd1305, 32'sd891, 32'sd547, 32'sd736, 32'sd930, 32'sd1600,
32'sd1289, 32'sd395, 32'sd912, 32'sd1049, 32'sd808, 32'sd420,
32'sd366, 32'sd1399, 32'sd357, 32'sd1222, 32'sd895, 32'sd310,
32'sd1314, 32'sd858, 32'sd1484, 32'sd1634, 32'sd1365, 32'sd1650,
32'sd1541, 32'sd181, 32'sd1159, 32'sd647, 32'sd510, 32'sd247,
32'sd295, 32'sd459, 32'sd250, 32'sd642, 32'sd1134, 32'sd1811,
32'sd1772, 32'sd892, 32'sd859, 32'sd115, 32'sd209, 32'sd1050,
32'sd792, 32'sd997, 32'sd343, 32'sd1695, 32'sd474, 32'sd1178,
32'sd233, 32'sd364, 32'sd855, 32'sd663, 32'sd1679, 32'sd889,
32'sd1046, 32'sd633, 32'sd963, 32'sd1638, 32'sd1945, 32'sd563,
32'sd787, 32'sd760, 32'sd1460, 32'sd1994, 32'sd1495, 32'sd216,
32'sd1365, 32'sd1936, 32'sd1218, 32'sd1100, 32'sd1979, 32'sd339,
32'sd272, 32'sd558, 32'sd570, 32'sd1734, 32'sd860, 32'sd1683,
32'sd1194, 32'sd1283, 32'sd446, 32'sd1991, 32'sd684, 32'sd1172,
32'sd387, 32'sd717, 32'sd1035, 32'sd1231, 32'sd975, 32'sd230,
32'sd1312, 32'sd1210, 32'sd888, 32'sd746, 32'sd1540, 32'sd492,
32'sd1205, 32'sd1011, 32'sd969, 32'sd1102, 32'sd1464, 32'sd401,
32'sd1478, 32'sd1391, 32'sd187, 32'sd1096, 32'sd203, 32'sd760,
32'sd1868, 32'sd1327, 32'sd413, 32'sd495, 32'sd162, 32'sd422,
32'sd1927, 32'sd890, 32'sd1050, 32'sd922, 32'sd138, 32'sd1438,
32'sd1128, 32'sd930, 32'sd1418, 32'sd1509, 32'sd1946, 32'sd1491,
32'sd664, 32'sd1842, 32'sd236, 32'sd1842, 32'sd1656, 32'sd1370,
32'sd1237, 32'sd1468, 32'sd1728, 32'sd840, 32'sd1144, 32'sd695,
32'sd1468, 32'sd401, 32'sd1730, 32'sd389, 32'sd1100, 32'sd874,
32'sd907, 32'sd1447, 32'sd649, 32'sd818, 32'sd1017, 32'sd1629,
32'sd289, 32'sd287, 32'sd843, 32'sd1287, 32'sd382, 32'sd1874,
32'sd173, 32'sd954, 32'sd384, 32'sd1493, 32'sd615, 32'sd1387,
32'sd744, 32'sd1224, 32'sd1014, 32'sd1265, 32'sd920, 32'sd1001,
32'sd620, 32'sd278, 32'sd1881, 32'sd1268, 32'sd1850, 32'sd555,
32'sd1773, 32'sd109, 32'sd287, 32'sd577, 32'sd981, 32'sd715,
32'sd1115, 32'sd1829, 32'sd181, 32'sd1470, 32'sd1131, 32'sd590,
32'sd884, 32'sd1108, 32'sd863, 32'sd1399, 32'sd805, 32'sd1669,
32'sd820, 32'sd1024, 32'sd1876, 32'sd1898, 32'sd1251, 32'sd215,
32'sd351, 32'sd1618, 32'sd1545, 32'sd1807, 32'sd858, 32'sd1594,
32'sd1411, 32'sd1722, 32'sd1685, 32'sd1934, 32'sd392, 32'sd171,
32'sd239, 32'sd154, 32'sd479, 32'sd1440, 32'sd405, 32'sd186,
32'sd976, 32'sd434, 32'sd1819, 32'sd1073, 32'sd1173, 32'sd741,
32'sd1718, 32'sd1229, 32'sd528, 32'sd740, 32'sd1627, 32'sd1451,
32'sd257, 32'sd217, 32'sd764, 32'sd445, 32'sd510, 32'sd516,
32'sd1888, 32'sd1630, 32'sd1110, 32'sd1746, 32'sd921, 32'sd1033,
32'sd449, 32'sd1975, 32'sd1317, 32'sd224, 32'sd1258, 32'sd1890,
32'sd488, 32'sd1384, 32'sd821, 32'sd1236, 32'sd1541, 32'sd146,
32'sd1416, 32'sd179, 32'sd1655, 32'sd656, 32'sd1734, 32'sd435,
32'sd870, 32'sd748, 32'sd1277, 32'sd194, 32'sd1529, 32'sd527,
32'sd617, 32'sd102, 32'sd1987, 32'sd1162, 32'sd1654, 32'sd906,
32'sd1348, 32'sd264, 32'sd1584, 32'sd1509, 32'sd1090, 32'sd244,
32'sd320, 32'sd1456, 32'sd486, 32'sd1358, 32'sd477, 32'sd890,
32'sd1364, 32'sd891, 32'sd173, 32'sd1735, 32'sd1280, 32'sd1730,
32'sd1828, 32'sd737, 32'sd927, 32'sd1189, 32'sd1266, 32'sd1202,
32'sd664, 32'sd1150, 32'sd1984, 32'sd1760, 32'sd1264, 32'sd426,
32'sd1660, 32'sd1529, 32'sd656, 32'sd1293, 32'sd1330, 32'sd264,
32'sd750, 32'sd1582, 32'sd1313, 32'sd235, 32'sd1060, 32'sd1789,
32'sd872, 32'sd827, 32'sd996, 32'sd1661, 32'sd1185, 32'sd622,
32'sd926, 32'sd1084, 32'sd1468, 32'sd208, 32'sd1092, 32'sd1535,
32'sd123, 32'sd1805, 32'sd1833, 32'sd779, 32'sd1459, 32'sd979,
32'sd803, 32'sd920, 32'sd1798, 32'sd142, 32'sd1449, 32'sd1598,
32'sd812, 32'sd990, 32'sd1526, 32'sd517, 32'sd417, 32'sd443,
32'sd1968, 32'sd110, 32'sd1225, 32'sd957, 32'sd1712, 32'sd1276,
32'sd676, 32'sd1266, 32'sd1573, 32'sd598, 32'sd251, 32'sd1753,
32'sd1228, 32'sd1165, 32'sd1843, 32'sd1785, 32'sd1807, 32'sd194,
32'sd416, 32'sd1310, 32'sd1700, 32'sd875, 32'sd1105, 32'sd1905,
32'sd1646, 32'sd1516, 32'sd1429, 32'sd328, 32'sd1399, 32'sd964,
32'sd1802, 32'sd1108, 32'sd196, 32'sd894, 32'sd1059, 32'sd1627,
32'sd533, 32'sd1601, 32'sd693, 32'sd1632, 32'sd1584, 32'sd391,
32'sd218, 32'sd879, 32'sd1386, 32'sd1089, 32'sd1447, 32'sd1999,
32'sd1763, 32'sd1402, 32'sd1929, 32'sd195, 32'sd628, 32'sd1256,
32'sd931, 32'sd1671, 32'sd812, 32'sd646, 32'sd194, 32'sd798,
32'sd1526, 32'sd1331, 32'sd1658, 32'sd1317, 32'sd1587, 32'sd164,
32'sd243, 32'sd1650, 32'sd1739, 32'sd597, 32'sd746, 32'sd1375,
32'sd1813, 32'sd1467, 32'sd198, 32'sd784, 32'sd176, 32'sd423,
32'sd669, 32'sd378, 32'sd192, 32'sd1455, 32'sd146, 32'sd1083,
32'sd1923, 32'sd1516, 32'sd1481, 32'sd1666, 32'sd1005, 32'sd328,
32'sd1024, 32'sd1179, 32'sd1686, 32'sd183, 32'sd985, 32'sd1845,
32'sd1669, 32'sd427, 32'sd286, 32'sd402, 32'sd126, 32'sd1218,
32'sd520, 32'sd1797, 32'sd673, 32'sd557, 32'sd1897, 32'sd1482,
32'sd1600, 32'sd1176, 32'sd768, 32'sd878, 32'sd1190, 32'sd620,
32'sd1357, 32'sd1295, 32'sd1320, 32'sd1104, 32'sd285, 32'sd728,
32'sd234, 32'sd649, 32'sd994, 32'sd1739, 32'sd639, 32'sd153,
32'sd1058, 32'sd152, 32'sd1307, 32'sd1401, 32'sd1133, 32'sd614,
32'sd617, 32'sd1470, 32'sd1661, 32'sd1427, 32'sd358, 32'sd420,
32'sd1539, 32'sd789, 32'sd1553, 32'sd1605, 32'sd1259, 32'sd1174,
32'sd650, 32'sd1667, 32'sd550, 32'sd715, 32'sd1273, 32'sd1359,
32'sd1777, 32'sd1613, 32'sd638, 32'sd133, 32'sd652, 32'sd1809,
32'sd357, 32'sd689, 32'sd1846, 32'sd1118, 32'sd1347, 32'sd899,
32'sd637, 32'sd700, 32'sd154, 32'sd1904, 32'sd1086, 32'sd1294,
32'sd670, 32'sd1390, 32'sd150, 32'sd1988, 32'sd633, 32'sd843,
32'sd945, 32'sd778, 32'sd987, 32'sd1643, 32'sd1797, 32'sd980,
32'sd1175, 32'sd1311, 32'sd1305, 32'sd1160, 32'sd789, 32'sd767,
32'sd131, 32'sd1349, 32'sd1428, 32'sd1621, 32'sd1419, 32'sd1988,
32'sd135, 32'sd706, 32'sd248, 32'sd1614, 32'sd563, 32'sd224,
32'sd182, 32'sd1524, 32'sd1778, 32'sd1089, 32'sd1403, 32'sd1706,
32'sd117, 32'sd590, 32'sd272, 32'sd746, 32'sd618, 32'sd1833,
32'sd1972, 32'sd1253, 32'sd1848, 32'sd1224, 32'sd647, 32'sd621,
32'sd1215, 32'sd1991, 32'sd1022, 32'sd362, 32'sd1846, 32'sd1649,
32'sd1785, 32'sd462, 32'sd1480, 32'sd1009, 32'sd1865, 32'sd558,
32'sd1281, 32'sd1868, 32'sd1444, 32'sd248, 32'sd1074, 32'sd1149,
32'sd1476, 32'sd1668, 32'sd660, 32'sd1603, 32'sd804, 32'sd137,
32'sd1603, 32'sd1860, 32'sd1190, 32'sd1675, 32'sd619, 32'sd855,
32'sd280, 32'sd1003, 32'sd258, 32'sd1081, 32'sd1486, 32'sd628,
32'sd1004, 32'sd883, 32'sd204, 32'sd934, 32'sd832, 32'sd509,
32'sd1410, 32'sd1665, 32'sd1220, 32'sd1985, 32'sd445, 32'sd1408,
32'sd916, 32'sd1730, 32'sd386, 32'sd539, 32'sd401, 32'sd1273,
32'sd1445, 32'sd1461, 32'sd684, 32'sd914, 32'sd927, 32'sd506,
32'sd1906, 32'sd372, 32'sd1249, 32'sd519, 32'sd666, 32'sd1498,
32'sd813, 32'sd1805, 32'sd164, 32'sd1131, 32'sd1259, 32'sd1054,
32'sd742, 32'sd238, 32'sd1578, 32'sd470, 32'sd1851, 32'sd1817,
32'sd1080, 32'sd575, 32'sd888, 32'sd719, 32'sd874, 32'sd1255,
32'sd1836, 32'sd1843, 32'sd874, 32'sd664, 32'sd947, 32'sd867,
32'sd1226, 32'sd294, 32'sd440, 32'sd1167, 32'sd1304, 32'sd1501,
32'sd1389, 32'sd1791, 32'sd1601, 32'sd875, 32'sd1298, 32'sd1914,
32'sd1537, 32'sd1752, 32'sd784, 32'sd1093, 32'sd1852, 32'sd880,
32'sd1174, 32'sd1080, 32'sd1088, 32'sd465, 32'sd891, 32'sd1216,
32'sd1989, 32'sd1079, 32'sd102, 32'sd739, 32'sd1158, 32'sd820,
32'sd706, 32'sd571, 32'sd1890, 32'sd745, 32'sd1379, 32'sd630,
32'sd1729, 32'sd1315, 32'sd1915, 32'sd525, 32'sd1034, 32'sd1681,
32'sd316, 32'sd1670, 32'sd1730, 32'sd1396, 32'sd143, 32'sd1976,
32'sd1518, 32'sd856, 32'sd446, 32'sd875, 32'sd828, 32'sd1899,
32'sd1773, 32'sd1581, 32'sd1217, 32'sd1310, 32'sd1363, 32'sd1781,
32'sd1870, 32'sd1495, 32'sd669, 32'sd979, 32'sd1664, 32'sd766,
32'sd746, 32'sd1699, 32'sd284, 32'sd133, 32'sd1961, 32'sd864,
32'sd953, 32'sd907, 32'sd736, 32'sd1989, 32'sd1370, 32'sd735,
32'sd966, 32'sd996, 32'sd946, 32'sd405, 32'sd801, 32'sd543,
32'sd674, 32'sd354, 32'sd1529, 32'sd485, 32'sd559, 32'sd1671,
32'sd913, 32'sd1922, 32'sd1226, 32'sd1715, 32'sd235, 32'sd1868,
32'sd1341, 32'sd989, 32'sd1291, 32'sd1417, 32'sd690, 32'sd772,
32'sd151, 32'sd951, 32'sd647, 32'sd1340, 32'sd852, 32'sd286,
32'sd1008, 32'sd1435, 32'sd1449, 32'sd510, 32'sd930, 32'sd739,
32'sd1862, 32'sd1025, 32'sd217, 32'sd731, 32'sd1155, 32'sd664,
32'sd1940, 32'sd188, 32'sd1063, 32'sd1621, 32'sd1862, 32'sd1140,
32'sd1947, 32'sd1195, 32'sd574, 32'sd237, 32'sd927, 32'sd1378,
32'sd1615, 32'sd1449, 32'sd315, 32'sd596, 32'sd1791, 32'sd243,
32'sd909, 32'sd801, 32'sd1698, 32'sd1037, 32'sd221, 32'sd1186,
32'sd1285, 32'sd153, 32'sd575, 32'sd1894, 32'sd1520, 32'sd751,
32'sd1343, 32'sd1449, 32'sd1851, 32'sd1276, 32'sd1866, 32'sd858,
32'sd1536, 32'sd1136, 32'sd1156, 32'sd225, 32'sd451, 32'sd1280,
32'sd1264, 32'sd501, 32'sd575, 32'sd920, 32'sd1264, 32'sd1781,
32'sd409, 32'sd1116, 32'sd1197, 32'sd1339, 32'sd1081, 32'sd887,
32'sd1349, 32'sd138, 32'sd880, 32'sd834, 32'sd726, 32'sd992,
32'sd1048, 32'sd566, 32'sd1751, 32'sd886, 32'sd1902, 32'sd1684,
32'sd597, 32'sd150, 32'sd181, 32'sd459, 32'sd1923, 32'sd568,
32'sd708, 32'sd1631, 32'sd347, 32'sd1261, 32'sd1052, 32'sd1939,
32'sd725, 32'sd1519, 32'sd448, 32'sd726, 32'sd1527, 32'sd703,
32'sd1285, 32'sd1823, 32'sd574, 32'sd686, 32'sd1142, 32'sd377,
32'sd1381, 32'sd1946, 32'sd140, 32'sd1336, 32'sd1730, 32'sd1502,
32'sd312, 32'sd1157, 32'sd151, 32'sd497, 32'sd761, 32'sd1654,
32'sd1808, 32'sd1437, 32'sd975, 32'sd101, 32'sd835, 32'sd687,
32'sd571, 32'sd347, 32'sd1092, 32'sd1488, 32'sd608, 32'sd1535,
32'sd660, 32'sd1382, 32'sd671, 32'sd1937, 32'sd263, 32'sd1833,
32'sd1222, 32'sd1438, 32'sd1336, 32'sd416, 32'sd942, 32'sd1936,
32'sd348, 32'sd825, 32'sd1035, 32'sd298, 32'sd627, 32'sd850,
32'sd278, 32'sd1498, 32'sd1074, 32'sd1119, 32'sd1065, 32'sd1229,
32'sd703, 32'sd1677, 32'sd479, 32'sd1918, 32'sd1281, 32'sd1826,
32'sd1612, 32'sd1114, 32'sd1443, 32'sd172, 32'sd893, 32'sd1211,
32'sd247, 32'sd356, 32'sd541, 32'sd255, 32'sd1513, 32'sd789,
32'sd1263, 32'sd569, 32'sd386, 32'sd1718, 32'sd509, 32'sd416,
32'sd749, 32'sd1707, 32'sd918, 32'sd1537, 32'sd688, 32'sd100,
32'sd437, 32'sd258, 32'sd350, 32'sd1292, 32'sd1531, 32'sd839,
32'sd1223, 32'sd685, 32'sd458, 32'sd813, 32'sd696, 32'sd1599,
32'sd1343, 32'sd700, 32'sd604, 32'sd1702, 32'sd631, 32'sd1732,
32'sd1233, 32'sd717, 32'sd1244, 32'sd1693, 32'sd1331, 32'sd263,
32'sd330, 32'sd993, 32'sd1207, 32'sd1639, 32'sd1936, 32'sd1221,
32'sd439, 32'sd1736, 32'sd950, 32'sd1546, 32'sd1863, 32'sd1056,
32'sd1962, 32'sd461, 32'sd389, 32'sd191, 32'sd1226, 32'sd622,
32'sd374, 32'sd1106, 32'sd1195, 32'sd1628, 32'sd387, 32'sd1722,
32'sd1022, 32'sd1142, 32'sd336, 32'sd1535, 32'sd1979, 32'sd393,
32'sd994, 32'sd1222, 32'sd1696, 32'sd907, 32'sd1217, 32'sd1043,
32'sd933, 32'sd444, 32'sd630, 32'sd1263, 32'sd617, 32'sd577,
32'sd895, 32'sd848, 32'sd890, 32'sd1844, 32'sd1597, 32'sd609,
32'sd1529, 32'sd1507, 32'sd1230, 32'sd1237, 32'sd396, 32'sd1533,
32'sd1085, 32'sd1890, 32'sd1892, 32'sd489, 32'sd773, 32'sd854,
32'sd1940, 32'sd1592, 32'sd1765, 32'sd1683, 32'sd473, 32'sd1805,
32'sd1636, 32'sd1673, 32'sd250, 32'sd1580, 32'sd1120, 32'sd443,
32'sd118, 32'sd860, 32'sd1651, 32'sd1657, 32'sd154, 32'sd780,
32'sd333, 32'sd1112, 32'sd1214, 32'sd669, 32'sd1856, 32'sd491,
32'sd830, 32'sd675, 32'sd225, 32'sd1588, 32'sd775, 32'sd1478,
32'sd978, 32'sd674, 32'sd409, 32'sd1614, 32'sd1354, 32'sd1632,
32'sd1784, 32'sd195, 32'sd896, 32'sd1556, 32'sd1182, 32'sd693,
32'sd349, 32'sd685, 32'sd998, 32'sd1832, 32'sd104, 32'sd184,
32'sd1105, 32'sd741, 32'sd1241, 32'sd1167, 32'sd308, 32'sd1903,
32'sd440, 32'sd1798, 32'sd904, 32'sd222, 32'sd236, 32'sd376,
32'sd405, 32'sd1961, 32'sd1084, 32'sd549, 32'sd385, 32'sd1595,
32'sd767, 32'sd844, 32'sd600, 32'sd132, 32'sd1441, 32'sd788,
32'sd278, 32'sd1951, 32'sd872, 32'sd1707, 32'sd109, 32'sd1773,
32'sd405, 32'sd1577, 32'sd447, 32'sd1752, 32'sd1972, 32'sd776,
32'sd739, 32'sd697, 32'sd1636, 32'sd1795, 32'sd527, 32'sd1255,
32'sd1317, 32'sd348, 32'sd523, 32'sd1025, 32'sd616, 32'sd1022,
32'sd1462, 32'sd1537, 32'sd739, 32'sd447, 32'sd1928, 32'sd483,
32'sd1280, 32'sd744, 32'sd1410, 32'sd907, 32'sd1717, 32'sd1216,
32'sd149, 32'sd681, 32'sd1800, 32'sd708, 32'sd1109, 32'sd1873,
32'sd436, 32'sd1827, 32'sd1178, 32'sd197, 32'sd1076, 32'sd674,
32'sd1201, 32'sd1584, 32'sd1326, 32'sd157, 32'sd269, 32'sd1817,
32'sd1696, 32'sd1897, 32'sd142, 32'sd365, 32'sd1141, 32'sd1153,
32'sd1678, 32'sd1163, 32'sd801, 32'sd1264, 32'sd1860, 32'sd897,
32'sd569, 32'sd351, 32'sd1011, 32'sd749, 32'sd1097, 32'sd731,
32'sd762, 32'sd173, 32'sd1769, 32'sd808, 32'sd115, 32'sd1673,
32'sd1871, 32'sd1960, 32'sd636, 32'sd1271, 32'sd326, 32'sd410,
32'sd1652, 32'sd1802, 32'sd756, 32'sd667, 32'sd704, 32'sd1000,
32'sd411, 32'sd1396, 32'sd475, 32'sd1405, 32'sd1043, 32'sd1716,
32'sd1480, 32'sd1520, 32'sd1001, 32'sd545, 32'sd1059, 32'sd195,
32'sd1976, 32'sd1865, 32'sd1556, 32'sd1868, 32'sd1333, 32'sd534,
32'sd459, 32'sd455, 32'sd1180, 32'sd268, 32'sd932, 32'sd141,
32'sd395, 32'sd1150, 32'sd1033, 32'sd1294, 32'sd674, 32'sd688,
32'sd447, 32'sd887, 32'sd516, 32'sd1877, 32'sd1834, 32'sd1816,
32'sd367, 32'sd896, 32'sd1173, 32'sd694, 32'sd1336, 32'sd1283,
32'sd832, 32'sd893, 32'sd644, 32'sd1775, 32'sd1022, 32'sd1693,
32'sd1408, 32'sd1657, 32'sd656, 32'sd733, 32'sd1618, 32'sd1651,
32'sd496, 32'sd884, 32'sd310, 32'sd811, 32'sd1873, 32'sd1463,
32'sd683, 32'sd1405, 32'sd1011, 32'sd1163, 32'sd633, 32'sd1019,
32'sd144, 32'sd593, 32'sd475, 32'sd1917, 32'sd1772, 32'sd1836,
32'sd1965, 32'sd904, 32'sd786, 32'sd1196, 32'sd107, 32'sd280,
32'sd932, 32'sd637, 32'sd1298, 32'sd401, 32'sd229, 32'sd655,
32'sd894, 32'sd1114, 32'sd1178, 32'sd737, 32'sd697, 32'sd1118,
32'sd162, 32'sd572, 32'sd674, 32'sd480, 32'sd1069, 32'sd1374,
32'sd1644, 32'sd1609, 32'sd348, 32'sd1724, 32'sd415, 32'sd661,
32'sd1090, 32'sd1000, 32'sd1723, 32'sd613, 32'sd1174, 32'sd162,
32'sd712, 32'sd349, 32'sd1286, 32'sd798, 32'sd1471, 32'sd1960,
32'sd921, 32'sd265, 32'sd1824, 32'sd919, 32'sd1517, 32'sd1831,
32'sd871, 32'sd1301, 32'sd1597, 32'sd1874, 32'sd714, 32'sd1404,
32'sd463, 32'sd480, 32'sd179, 32'sd1554, 32'sd1742, 32'sd517,
32'sd774, 32'sd535, 32'sd134, 32'sd1106, 32'sd378, 32'sd1959,
32'sd1829, 32'sd1834, 32'sd1709, 32'sd286, 32'sd1573, 32'sd1345,
32'sd1509, 32'sd1744, 32'sd1751, 32'sd416, 32'sd1767, 32'sd699,
32'sd233, 32'sd1574, 32'sd1684, 32'sd1823, 32'sd1301, 32'sd1125,
32'sd116, 32'sd132, 32'sd608, 32'sd358, 32'sd1379, 32'sd719,
32'sd510, 32'sd1605, 32'sd1265, 32'sd900, 32'sd380, 32'sd1921,
32'sd445, 32'sd1159, 32'sd1901, 32'sd1168, 32'sd823, 32'sd1850,
32'sd430, 32'sd1627, 32'sd1306, 32'sd1791, 32'sd131, 32'sd601,
32'sd971, 32'sd758, 32'sd547, 32'sd1233, 32'sd1524, 32'sd1898,
32'sd1158, 32'sd1922, 32'sd564, 32'sd1369, 32'sd1343, 32'sd1700,
32'sd1371, 32'sd1026, 32'sd1388, 32'sd647, 32'sd1317, 32'sd1565,
32'sd1884, 32'sd554, 32'sd601, 32'sd1217, 32'sd1926, 32'sd1618,
32'sd1057, 32'sd1317, 32'sd1270, 32'sd371, 32'sd1536, 32'sd1980,
32'sd877, 32'sd322, 32'sd607, 32'sd392, 32'sd888, 32'sd657,
32'sd272, 32'sd1947, 32'sd337, 32'sd476, 32'sd1966, 32'sd1658,
32'sd875, 32'sd959, 32'sd1967, 32'sd168, 32'sd1771, 32'sd1968,
32'sd641, 32'sd1568, 32'sd1663, 32'sd450, 32'sd1960, 32'sd1594,
32'sd572, 32'sd191, 32'sd595, 32'sd1007, 32'sd1091, 32'sd768,
32'sd1427, 32'sd111, 32'sd1586, 32'sd1061, 32'sd1369, 32'sd1141,
32'sd718, 32'sd388, 32'sd1591, 32'sd1502, 32'sd444, 32'sd984,
32'sd1157, 32'sd1274, 32'sd864, 32'sd1875, 32'sd609, 32'sd224,
32'sd1652, 32'sd660, 32'sd543, 32'sd1463, 32'sd1446, 32'sd544,
32'sd186, 32'sd464, 32'sd1450, 32'sd942, 32'sd1520, 32'sd1868,
32'sd266, 32'sd1339, 32'sd963, 32'sd1521, 32'sd398, 32'sd1448,
32'sd382, 32'sd1179, 32'sd883, 32'sd786, 32'sd1574, 32'sd151,
32'sd225, 32'sd895, 32'sd1551, 32'sd1657, 32'sd1501, 32'sd274,
32'sd1909, 32'sd1773, 32'sd1707, 32'sd1284, 32'sd1950, 32'sd699,
32'sd1861, 32'sd322, 32'sd961, 32'sd838, 32'sd1089, 32'sd995,
32'sd703, 32'sd680, 32'sd1871, 32'sd1319, 32'sd236, 32'sd1667,
32'sd1468, 32'sd1142, 32'sd937, 32'sd426, 32'sd175, 32'sd800,
32'sd591, 32'sd1554, 32'sd127, 32'sd483, 32'sd1220, 32'sd1607,
32'sd272, 32'sd1241, 32'sd873, 32'sd625, 32'sd1719, 32'sd808,
32'sd1754, 32'sd1069, 32'sd798, 32'sd1344, 32'sd280, 32'sd1153,
32'sd441, 32'sd1994, 32'sd1474, 32'sd1074, 32'sd1412, 32'sd758,
32'sd1235, 32'sd1497, 32'sd1902, 32'sd1874, 32'sd1803, 32'sd1663,
32'sd1859, 32'sd1003, 32'sd1881, 32'sd1681, 32'sd103, 32'sd843,
32'sd1866, 32'sd1458, 32'sd1766, 32'sd1401, 32'sd781, 32'sd1888,
32'sd1854, 32'sd1459, 32'sd1742, 32'sd625, 32'sd103, 32'sd311,
32'sd1325, 32'sd173, 32'sd1446, 32'sd1296, 32'sd1259, 32'sd374,
32'sd763, 32'sd130, 32'sd648, 32'sd1112, 32'sd651, 32'sd1782,
32'sd103, 32'sd1014, 32'sd973, 32'sd121, 32'sd442, 32'sd999,
32'sd356, 32'sd1269, 32'sd1774, 32'sd1032, 32'sd440, 32'sd447,
32'sd1496, 32'sd1203, 32'sd199, 32'sd1659, 32'sd921, 32'sd886,
32'sd504, 32'sd498, 32'sd261, 32'sd1613, 32'sd608, 32'sd1969,
32'sd513, 32'sd1121, 32'sd1342, 32'sd1893, 32'sd1860, 32'sd1915,
32'sd1149, 32'sd635, 32'sd1895, 32'sd1077, 32'sd1974, 32'sd153,
32'sd1283, 32'sd1030, 32'sd651, 32'sd808, 32'sd1971, 32'sd1296,
32'sd1177, 32'sd1942, 32'sd731, 32'sd1954, 32'sd835, 32'sd1391,
32'sd1766, 32'sd1256, 32'sd291, 32'sd106, 32'sd952, 32'sd1781,
32'sd1405, 32'sd1340, 32'sd520, 32'sd532, 32'sd652, 32'sd809,
32'sd1833, 32'sd423, 32'sd1371, 32'sd1057, 32'sd363, 32'sd1613,
32'sd326, 32'sd1140, 32'sd848, 32'sd299, 32'sd807, 32'sd1487,
32'sd349, 32'sd382, 32'sd364, 32'sd1037, 32'sd879, 32'sd1102,
32'sd1446, 32'sd299, 32'sd1323, 32'sd402, 32'sd1218, 32'sd1400,
32'sd595, 32'sd1032, 32'sd216, 32'sd1072, 32'sd1881, 32'sd1947,
32'sd1778, 32'sd350, 32'sd1460, 32'sd859, 32'sd1009, 32'sd323,
32'sd1732, 32'sd555, 32'sd1871, 32'sd395, 32'sd1206, 32'sd1107,
32'sd174, 32'sd1217, 32'sd261, 32'sd1638, 32'sd1605, 32'sd472,
32'sd822, 32'sd712, 32'sd1310, 32'sd1896, 32'sd1536, 32'sd944,
32'sd195, 32'sd1856, 32'sd1361, 32'sd1487, 32'sd1624, 32'sd1482,
32'sd469, 32'sd985, 32'sd1723, 32'sd1287, 32'sd1704, 32'sd1689,
32'sd1812, 32'sd1679, 32'sd252, 32'sd550, 32'sd510, 32'sd528,
32'sd1092, 32'sd1452, 32'sd878, 32'sd823, 32'sd706, 32'sd362,
32'sd790, 32'sd834, 32'sd864, 32'sd823, 32'sd976, 32'sd1843,
32'sd663, 32'sd1799, 32'sd192, 32'sd403, 32'sd270, 32'sd1695,
32'sd1304, 32'sd1434, 32'sd535, 32'sd1641, 32'sd1317, 32'sd1698,
32'sd944, 32'sd1668, 32'sd1096, 32'sd1372, 32'sd792, 32'sd1766,
32'sd1971, 32'sd712, 32'sd1731, 32'sd1296, 32'sd648, 32'sd169,
32'sd838, 32'sd592, 32'sd1253, 32'sd1733, 32'sd720, 32'sd661,
32'sd827, 32'sd1828, 32'sd1935, 32'sd240, 32'sd185, 32'sd273,
32'sd1777, 32'sd1471, 32'sd1054, 32'sd483, 32'sd841, 32'sd1079,
32'sd693, 32'sd1774, 32'sd526, 32'sd1039, 32'sd1712, 32'sd368,
32'sd892, 32'sd1404, 32'sd184, 32'sd1893, 32'sd1622, 32'sd1233,
32'sd1945, 32'sd479, 32'sd567, 32'sd362, 32'sd1743, 32'sd1889,
32'sd817, 32'sd866, 32'sd718, 32'sd782, 32'sd1380, 32'sd250,
32'sd1322, 32'sd1301, 32'sd1055, 32'sd1214, 32'sd279, 32'sd1079,
32'sd1275, 32'sd1343, 32'sd1809, 32'sd374, 32'sd1273, 32'sd264,
32'sd1182, 32'sd355, 32'sd1220, 32'sd1089, 32'sd427, 32'sd616,
32'sd527, 32'sd427, 32'sd281, 32'sd1668, 32'sd126, 32'sd517,
32'sd1284, 32'sd685, 32'sd339, 32'sd1370, 32'sd589, 32'sd1584,
32'sd1440, 32'sd1508, 32'sd520, 32'sd870, 32'sd1284, 32'sd298,
32'sd369, 32'sd778, 32'sd1415, 32'sd945, 32'sd535, 32'sd295,
32'sd1630, 32'sd843, 32'sd1641, 32'sd1992, 32'sd715, 32'sd559,
32'sd1057, 32'sd1167, 32'sd1533, 32'sd1452, 32'sd848, 32'sd375,
32'sd1679, 32'sd167, 32'sd164, 32'sd1270, 32'sd1223, 32'sd909,
32'sd204, 32'sd553, 32'sd1611, 32'sd1647, 32'sd1762, 32'sd1230,
32'sd1675, 32'sd1014, 32'sd200, 32'sd1409, 32'sd210, 32'sd944,
32'sd1642, 32'sd1639, 32'sd1162, 32'sd1472, 32'sd1275, 32'sd1582,
32'sd402, 32'sd1151, 32'sd970, 32'sd1963, 32'sd1220, 32'sd1031,
32'sd1321, 32'sd897, 32'sd1123, 32'sd1221, 32'sd908, 32'sd338,
32'sd536, 32'sd1170, 32'sd364, 32'sd1287, 32'sd1960, 32'sd578,
32'sd1354, 32'sd936, 32'sd1786, 32'sd699, 32'sd1863, 32'sd1345,
32'sd538, 32'sd715, 32'sd205, 32'sd405, 32'sd601, 32'sd1490,
32'sd1391, 32'sd1979, 32'sd1676, 32'sd860, 32'sd646, 32'sd1224,
32'sd1413, 32'sd965, 32'sd1612, 32'sd1122, 32'sd684, 32'sd1647,
32'sd148, 32'sd838, 32'sd1776, 32'sd559, 32'sd1717, 32'sd1265,
32'sd1742, 32'sd226, 32'sd168, 32'sd100, 32'sd1934, 32'sd259,
32'sd1896, 32'sd774, 32'sd1233, 32'sd1865, 32'sd1537, 32'sd1034,
32'sd1045, 32'sd764, 32'sd998, 32'sd1194, 32'sd1404, 32'sd1761,
32'sd687, 32'sd1496, 32'sd842, 32'sd1448, 32'sd636, 32'sd1231,
32'sd694, 32'sd1691, 32'sd1376, 32'sd204, 32'sd1365, 32'sd677,
32'sd949, 32'sd1583, 32'sd959, 32'sd1551, 32'sd238, 32'sd1677,
32'sd1019, 32'sd728, 32'sd1987, 32'sd386, 32'sd1524, 32'sd716,
32'sd790, 32'sd1979, 32'sd305, 32'sd445, 32'sd1218, 32'sd833,
32'sd643, 32'sd1424, 32'sd895, 32'sd192, 32'sd149, 32'sd365,
32'sd2000, 32'sd1345, 32'sd862, 32'sd859, 32'sd1250, 32'sd946,
32'sd455, 32'sd440, 32'sd847, 32'sd551, 32'sd435, 32'sd842,
32'sd117, 32'sd688, 32'sd402, 32'sd289, 32'sd1363, 32'sd1661,
32'sd693, 32'sd1257, 32'sd147, 32'sd1895, 32'sd839, 32'sd220,
32'sd191, 32'sd1706, 32'sd434, 32'sd215, 32'sd1439, 32'sd1565,
32'sd871, 32'sd1709, 32'sd825, 32'sd260, 32'sd1515, 32'sd440,
32'sd1543, 32'sd545, 32'sd1082, 32'sd1608, 32'sd746, 32'sd1444,
32'sd849, 32'sd1269, 32'sd169, 32'sd909, 32'sd691, 32'sd1966,
32'sd1940, 32'sd1276, 32'sd445, 32'sd993, 32'sd1421, 32'sd1545,
32'sd1274, 32'sd181, 32'sd266, 32'sd1538, 32'sd1924, 32'sd1315,
32'sd185, 32'sd207, 32'sd873, 32'sd1848, 32'sd165, 32'sd301,
32'sd1902, 32'sd853, 32'sd458, 32'sd1241, 32'sd891, 32'sd645,
32'sd1311, 32'sd998, 32'sd1309, 32'sd456, 32'sd137, 32'sd399,
32'sd230, 32'sd525, 32'sd689, 32'sd1161, 32'sd1456, 32'sd915,
32'sd757, 32'sd652, 32'sd480, 32'sd1782, 32'sd1847, 32'sd273,
32'sd1186, 32'sd629, 32'sd1786, 32'sd1565, 32'sd1470, 32'sd210,
32'sd457, 32'sd187, 32'sd716, 32'sd1302, 32'sd1254, 32'sd1479,
32'sd1911, 32'sd1435, 32'sd949, 32'sd504, 32'sd775, 32'sd1452,
32'sd1700, 32'sd1341, 32'sd1390, 32'sd1245, 32'sd449, 32'sd1503,
32'sd674, 32'sd1994, 32'sd704, 32'sd409, 32'sd432, 32'sd929,
32'sd1697, 32'sd1902, 32'sd1939, 32'sd506, 32'sd1717, 32'sd1637,
32'sd571, 32'sd820, 32'sd594, 32'sd1874, 32'sd1112, 32'sd513,
32'sd1761, 32'sd1445, 32'sd1912, 32'sd308, 32'sd433, 32'sd1765,
32'sd1473, 32'sd1549, 32'sd169, 32'sd1476, 32'sd1239, 32'sd1450,
32'sd1116, 32'sd1498, 32'sd445, 32'sd597, 32'sd312, 32'sd412,
32'sd1801, 32'sd1521, 32'sd1830, 32'sd1111, 32'sd529, 32'sd891,
32'sd868, 32'sd822, 32'sd1066, 32'sd543, 32'sd1351, 32'sd844,
32'sd785, 32'sd953, 32'sd981, 32'sd1101, 32'sd973, 32'sd1201,
32'sd1554, 32'sd1860, 32'sd481, 32'sd1204, 32'sd1157, 32'sd1537,
32'sd1793, 32'sd742, 32'sd1594, 32'sd1700, 32'sd1551, 32'sd1169,
32'sd1270, 32'sd1120, 32'sd1091, 32'sd1458, 32'sd1810, 32'sd692,
32'sd240, 32'sd1859, 32'sd351, 32'sd1338, 32'sd477, 32'sd633,
32'sd366, 32'sd995, 32'sd1176, 32'sd1247, 32'sd1271, 32'sd535,
32'sd1550, 32'sd207, 32'sd307, 32'sd470, 32'sd1107, 32'sd848,
32'sd1864, 32'sd1521, 32'sd385, 32'sd971, 32'sd468, 32'sd357,
32'sd900, 32'sd156, 32'sd1826, 32'sd464, 32'sd695, 32'sd622,
32'sd741, 32'sd206, 32'sd1930, 32'sd1694, 32'sd1165, 32'sd1339,
32'sd1725, 32'sd1454, 32'sd1551, 32'sd1131, 32'sd1721, 32'sd1645,
32'sd1802, 32'sd1328, 32'sd849, 32'sd1831, 32'sd292, 32'sd1384,
32'sd1576, 32'sd437, 32'sd253, 32'sd623, 32'sd1943, 32'sd1984,
32'sd1564, 32'sd999, 32'sd878, 32'sd1595, 32'sd1111, 32'sd1533,
32'sd603, 32'sd748, 32'sd1263, 32'sd1475, 32'sd1965, 32'sd1104,
32'sd1185, 32'sd652, 32'sd1895, 32'sd900, 32'sd334, 32'sd729,
32'sd1418, 32'sd1555, 32'sd529, 32'sd1182, 32'sd1788, 32'sd1902,
32'sd1588, 32'sd1396, 32'sd305, 32'sd1491, 32'sd1152, 32'sd1519,
32'sd912, 32'sd933, 32'sd1247, 32'sd918, 32'sd1347, 32'sd1784,
32'sd228, 32'sd493, 32'sd1203, 32'sd749, 32'sd1636, 32'sd413,
32'sd963, 32'sd1358, 32'sd1746, 32'sd854, 32'sd1121, 32'sd1581,
32'sd1939, 32'sd286, 32'sd828, 32'sd1826, 32'sd125, 32'sd1133,
32'sd1782, 32'sd1374, 32'sd439, 32'sd1767, 32'sd1520, 32'sd780,
32'sd516, 32'sd1598, 32'sd1731, 32'sd202, 32'sd1332, 32'sd1655,
32'sd783, 32'sd911, 32'sd879, 32'sd1079, 32'sd1933, 32'sd1814,
32'sd1306, 32'sd1003, 32'sd1144, 32'sd965, 32'sd383, 32'sd1222,
32'sd1755, 32'sd460, 32'sd1516, 32'sd1847, 32'sd995, 32'sd521,
32'sd866, 32'sd1398, 32'sd807, 32'sd1869, 32'sd1349, 32'sd1483,
32'sd1968, 32'sd982, 32'sd678, 32'sd1401, 32'sd613, 32'sd555,
32'sd645, 32'sd962, 32'sd1429, 32'sd1939, 32'sd572, 32'sd502,
32'sd658, 32'sd1298, 32'sd1924, 32'sd801, 32'sd1922, 32'sd542,
32'sd611, 32'sd1673, 32'sd721, 32'sd1734, 32'sd1737, 32'sd1590,
32'sd1532, 32'sd714, 32'sd1954, 32'sd848, 32'sd1434, 32'sd1955,
32'sd553, 32'sd848, 32'sd577, 32'sd1831, 32'sd809, 32'sd1529,
32'sd1953, 32'sd1720, 32'sd1504, 32'sd1493, 32'sd1442, 32'sd763,
32'sd329, 32'sd1228, 32'sd588, 32'sd1153, 32'sd670, 32'sd1144,
32'sd100, 32'sd1394, 32'sd1240, 32'sd802, 32'sd1837, 32'sd265,
32'sd614, 32'sd460, 32'sd1314, 32'sd1108, 32'sd527, 32'sd887,
32'sd1196, 32'sd1617, 32'sd532, 32'sd1239, 32'sd143, 32'sd855,
32'sd1176, 32'sd822, 32'sd1097, 32'sd590, 32'sd1130, 32'sd1171,
32'sd623, 32'sd1976, 32'sd1806, 32'sd1317, 32'sd1549, 32'sd672,
32'sd1119, 32'sd749, 32'sd534, 32'sd1675, 32'sd1990, 32'sd1934,
32'sd551, 32'sd131, 32'sd323, 32'sd1801, 32'sd1675, 32'sd1494,
32'sd1993, 32'sd1951, 32'sd425, 32'sd918, 32'sd781, 32'sd1202,
32'sd1024, 32'sd782, 32'sd697, 32'sd380, 32'sd1094, 32'sd535,
32'sd545, 32'sd706, 32'sd1852, 32'sd584, 32'sd1984, 32'sd687,
32'sd753, 32'sd1099, 32'sd1065, 32'sd1853, 32'sd1095, 32'sd1711,
32'sd1205, 32'sd1668, 32'sd1591, 32'sd1873, 32'sd979, 32'sd504,
32'sd243, 32'sd848, 32'sd590, 32'sd666, 32'sd1610, 32'sd247,
32'sd1228, 32'sd1518, 32'sd1869, 32'sd1545, 32'sd1493, 32'sd894,
32'sd462, 32'sd936, 32'sd1320, 32'sd892, 32'sd1707, 32'sd1368,
32'sd822, 32'sd541, 32'sd1646, 32'sd535, 32'sd502, 32'sd134,
32'sd1679, 32'sd1802, 32'sd1697, 32'sd1129, 32'sd468, 32'sd1614,
32'sd225, 32'sd153, 32'sd324, 32'sd1354, 32'sd1779, 32'sd1805,
32'sd379, 32'sd1903, 32'sd1269, 32'sd750, 32'sd410, 32'sd1506,
32'sd319, 32'sd1853, 32'sd206, 32'sd785, 32'sd1636, 32'sd1676,
32'sd1995, 32'sd983, 32'sd1209, 32'sd158, 32'sd1351, 32'sd1244,
32'sd1712, 32'sd849, 32'sd1086, 32'sd1591, 32'sd1150, 32'sd1861,
32'sd148, 32'sd1112, 32'sd830, 32'sd1241, 32'sd783, 32'sd655,
32'sd1317, 32'sd1814, 32'sd249, 32'sd1987, 32'sd699, 32'sd428,
32'sd776, 32'sd913, 32'sd1198, 32'sd363, 32'sd1415, 32'sd1882,
32'sd780, 32'sd633, 32'sd1575, 32'sd1900, 32'sd204, 32'sd1940,
32'sd1387, 32'sd309, 32'sd718, 32'sd1236, 32'sd1631, 32'sd1995,
32'sd1194, 32'sd1520, 32'sd288, 32'sd366, 32'sd1639, 32'sd1602,
32'sd840, 32'sd224, 32'sd986, 32'sd277, 32'sd494, 32'sd1975,
32'sd1328, 32'sd1911, 32'sd1985, 32'sd1261, 32'sd1733, 32'sd1607,
32'sd1247, 32'sd1304, 32'sd1809, 32'sd729, 32'sd153, 32'sd1164,
32'sd636, 32'sd1366, 32'sd778, 32'sd1296, 32'sd1610, 32'sd309,
32'sd760, 32'sd959, 32'sd1040, 32'sd375, 32'sd1217, 32'sd121,
32'sd1212, 32'sd1665, 32'sd613, 32'sd902, 32'sd960, 32'sd571,
32'sd1206, 32'sd1793, 32'sd275, 32'sd387, 32'sd256, 32'sd407,
32'sd1777, 32'sd752, 32'sd1857, 32'sd1828, 32'sd1366, 32'sd1817,
32'sd1197, 32'sd1492, 32'sd891, 32'sd455, 32'sd457, 32'sd1162,
32'sd114, 32'sd1455, 32'sd1383, 32'sd277, 32'sd1864, 32'sd204,
32'sd229, 32'sd485, 32'sd1156, 32'sd673, 32'sd970, 32'sd928,
32'sd930, 32'sd1444, 32'sd1817, 32'sd1105, 32'sd1845, 32'sd237,
32'sd1101, 32'sd1925, 32'sd1996, 32'sd909, 32'sd1640, 32'sd1273,
32'sd430, 32'sd1516, 32'sd1471, 32'sd1502, 32'sd1981, 32'sd204,
32'sd934, 32'sd175, 32'sd268, 32'sd1769, 32'sd499, 32'sd638,
32'sd1405, 32'sd1945, 32'sd1621, 32'sd447, 32'sd1625, 32'sd302,
32'sd193, 32'sd405, 32'sd333, 32'sd1018, 32'sd272, 32'sd148,
32'sd1333, 32'sd1513, 32'sd1358, 32'sd125, 32'sd1793, 32'sd1914,
32'sd131, 32'sd323, 32'sd533, 32'sd935, 32'sd1045, 32'sd318,
32'sd1331, 32'sd942, 32'sd1240, 32'sd573, 32'sd994, 32'sd660,
32'sd597, 32'sd1740, 32'sd266, 32'sd115, 32'sd1356, 32'sd271,
32'sd100, 32'sd1368, 32'sd317, 32'sd1840, 32'sd488, 32'sd1883,
32'sd1014, 32'sd1905, 32'sd1508, 32'sd615, 32'sd1774, 32'sd487,
32'sd929, 32'sd1893, 32'sd441, 32'sd244, 32'sd1504, 32'sd328,
32'sd1683, 32'sd462, 32'sd1362, 32'sd1827, 32'sd911, 32'sd614,
32'sd1544, 32'sd1641, 32'sd1673, 32'sd669, 32'sd1016, 32'sd389,
32'sd1239, 32'sd833, 32'sd395, 32'sd1421, 32'sd1292, 32'sd124,
32'sd1828, 32'sd1374, 32'sd864, 32'sd901, 32'sd1208, 32'sd463,
32'sd1202, 32'sd1634, 32'sd1150, 32'sd1733, 32'sd1068, 32'sd182,
32'sd1667, 32'sd1866, 32'sd1815, 32'sd1164, 32'sd350, 32'sd356,
32'sd1073, 32'sd1309, 32'sd1380, 32'sd220, 32'sd1603, 32'sd1109,
32'sd1677, 32'sd125, 32'sd1215, 32'sd819, 32'sd1615, 32'sd1041,
32'sd1068, 32'sd1489, 32'sd1342, 32'sd1179, 32'sd465, 32'sd1015,
32'sd260, 32'sd1115, 32'sd1916, 32'sd1930, 32'sd945, 32'sd1859,
32'sd348, 32'sd1573, 32'sd379, 32'sd1316, 32'sd1423, 32'sd1529,
32'sd1735, 32'sd356, 32'sd1113, 32'sd1568, 32'sd589, 32'sd1507,
32'sd722, 32'sd1822, 32'sd229, 32'sd146, 32'sd1810, 32'sd1497,
32'sd1413, 32'sd1515, 32'sd532, 32'sd350, 32'sd672, 32'sd662,
32'sd1202, 32'sd689, 32'sd1747, 32'sd1920, 32'sd1939, 32'sd1113,
32'sd1675, 32'sd441, 32'sd1712, 32'sd917, 32'sd813, 32'sd524,
32'sd771, 32'sd752, 32'sd1890, 32'sd1063, 32'sd1018, 32'sd1390,
32'sd1307, 32'sd1111, 32'sd1555, 32'sd246, 32'sd1604, 32'sd1645,
32'sd1412, 32'sd390, 32'sd1873, 32'sd224, 32'sd576, 32'sd1733,
32'sd1778, 32'sd377, 32'sd1978, 32'sd110, 32'sd1825, 32'sd1609,
32'sd1262, 32'sd1673, 32'sd461, 32'sd1657, 32'sd1538, 32'sd624,
32'sd414, 32'sd1462, 32'sd1050, 32'sd262, 32'sd411, 32'sd1489,
32'sd848, 32'sd315, 32'sd672, 32'sd147, 32'sd502, 32'sd1979,
32'sd416, 32'sd1483, 32'sd1630, 32'sd1499, 32'sd873, 32'sd1462,
32'sd912, 32'sd1356, 32'sd1080, 32'sd824, 32'sd251, 32'sd1650,
32'sd346, 32'sd741, 32'sd1566, 32'sd1796, 32'sd1717, 32'sd391,
32'sd1660, 32'sd600, 32'sd408, 32'sd1419, 32'sd108, 32'sd799,
32'sd1480, 32'sd926, 32'sd845, 32'sd724, 32'sd319, 32'sd1392,
32'sd830, 32'sd1237, 32'sd359, 32'sd843, 32'sd672, 32'sd1484,
32'sd186, 32'sd831, 32'sd1544, 32'sd998, 32'sd1374, 32'sd1814,
32'sd1668, 32'sd1365, 32'sd1724, 32'sd1467, 32'sd1501, 32'sd1869,
32'sd122, 32'sd1449, 32'sd122, 32'sd1687, 32'sd1150, 32'sd1965,
32'sd980, 32'sd489, 32'sd670, 32'sd697, 32'sd1987, 32'sd153,
32'sd1222, 32'sd1206, 32'sd1259, 32'sd1040, 32'sd869, 32'sd490,
32'sd1137, 32'sd814, 32'sd300, 32'sd1395, 32'sd1136, 32'sd828,
32'sd1073, 32'sd1455, 32'sd152, 32'sd1949, 32'sd615, 32'sd971,
32'sd731, 32'sd436, 32'sd1695, 32'sd101, 32'sd1329, 32'sd1691,
32'sd905, 32'sd960, 32'sd1305, 32'sd618, 32'sd1161, 32'sd1612,
32'sd856, 32'sd380, 32'sd376, 32'sd930, 32'sd223, 32'sd544,
32'sd1755, 32'sd864, 32'sd1488, 32'sd995, 32'sd466, 32'sd1185,
32'sd179, 32'sd242, 32'sd1223, 32'sd665, 32'sd215, 32'sd164,
32'sd440, 32'sd689, 32'sd1373, 32'sd1338, 32'sd424, 32'sd1929,
32'sd1346, 32'sd1186, 32'sd1118, 32'sd1597, 32'sd1814, 32'sd1663,
32'sd1034, 32'sd522, 32'sd1706, 32'sd815, 32'sd170, 32'sd1379,
32'sd1321, 32'sd1275, 32'sd1687, 32'sd1175, 32'sd1564, 32'sd489,
32'sd1889, 32'sd1122, 32'sd918, 32'sd141, 32'sd307, 32'sd931,
32'sd1566, 32'sd1707, 32'sd714, 32'sd284, 32'sd1331, 32'sd1926,
32'sd291, 32'sd1065, 32'sd1009, 32'sd498, 32'sd1236, 32'sd312,
32'sd1297, 32'sd913, 32'sd1328, 32'sd1133, 32'sd1686, 32'sd1297,
32'sd1782, 32'sd1561, 32'sd920, 32'sd1561, 32'sd242, 32'sd1735,
32'sd1440, 32'sd238, 32'sd1351, 32'sd1489, 32'sd1757, 32'sd716,
32'sd657, 32'sd192, 32'sd946, 32'sd1196, 32'sd401, 32'sd653,
32'sd1217, 32'sd780, 32'sd970, 32'sd1098, 32'sd1643, 32'sd526,
32'sd1085, 32'sd396, 32'sd867, 32'sd1767, 32'sd263, 32'sd1853,
32'sd875, 32'sd413, 32'sd1825, 32'sd1621, 32'sd930, 32'sd620,
32'sd1646, 32'sd1408, 32'sd1278, 32'sd1142, 32'sd924, 32'sd1423,
32'sd575, 32'sd1308, 32'sd737, 32'sd1902, 32'sd1725, 32'sd1798,
32'sd1151, 32'sd787, 32'sd623, 32'sd1624, 32'sd298, 32'sd808,
32'sd953, 32'sd855, 32'sd172, 32'sd666, 32'sd479, 32'sd376,
32'sd1834, 32'sd1477, 32'sd1282, 32'sd501, 32'sd659, 32'sd1430,
32'sd852, 32'sd1216, 32'sd1785, 32'sd1352, 32'sd389, 32'sd243,
32'sd1921, 32'sd1083, 32'sd1061, 32'sd139, 32'sd338, 32'sd1581,
32'sd752, 32'sd1965, 32'sd554, 32'sd1182, 32'sd729, 32'sd315,
32'sd483, 32'sd1832, 32'sd1716, 32'sd127, 32'sd703, 32'sd1259,
32'sd787, 32'sd1808, 32'sd959, 32'sd1386, 32'sd213, 32'sd384,
32'sd1380, 32'sd1905, 32'sd893, 32'sd1568, 32'sd1361, 32'sd1271,
32'sd1236, 32'sd1349, 32'sd143, 32'sd1387, 32'sd1725, 32'sd1540,
32'sd1180, 32'sd1545, 32'sd1831, 32'sd1659, 32'sd670, 32'sd103,
32'sd399, 32'sd1833, 32'sd212, 32'sd1981, 32'sd230, 32'sd807,
32'sd813, 32'sd680, 32'sd1509, 32'sd930, 32'sd745, 32'sd239,
32'sd603, 32'sd566, 32'sd1702, 32'sd128, 32'sd1008, 32'sd1161,
32'sd1739, 32'sd1194, 32'sd552, 32'sd747, 32'sd1071, 32'sd429,
32'sd1477, 32'sd426, 32'sd1743, 32'sd551, 32'sd1335, 32'sd1241,
32'sd1359, 32'sd165, 32'sd1415, 32'sd1870, 32'sd1083, 32'sd1395,
32'sd792, 32'sd1022, 32'sd612, 32'sd1125, 32'sd1548, 32'sd766,
32'sd1318, 32'sd1327, 32'sd1221, 32'sd1605, 32'sd1659, 32'sd1665,
32'sd871, 32'sd1726, 32'sd1103, 32'sd672, 32'sd628, 32'sd715,
32'sd1077, 32'sd716, 32'sd1394, 32'sd815, 32'sd1284, 32'sd1869,
32'sd1965, 32'sd1680, 32'sd1976, 32'sd1496, 32'sd1242, 32'sd730,
32'sd791, 32'sd675, 32'sd383, 32'sd604, 32'sd1225, 32'sd1446,
32'sd1647, 32'sd180, 32'sd346, 32'sd1345, 32'sd1443, 32'sd928,
32'sd622, 32'sd864, 32'sd157, 32'sd888, 32'sd1216, 32'sd1433,
32'sd652, 32'sd1804, 32'sd580, 32'sd807, 32'sd1891, 32'sd1725,
32'sd831, 32'sd610, 32'sd1070, 32'sd243, 32'sd1824, 32'sd1980,
32'sd159, 32'sd1732, 32'sd1891, 32'sd1567, 32'sd669, 32'sd1731,
32'sd254, 32'sd845, 32'sd1380, 32'sd857, 32'sd266, 32'sd1545,
32'sd183, 32'sd1423, 32'sd196, 32'sd925, 32'sd1958, 32'sd1773,
32'sd287, 32'sd173, 32'sd518, 32'sd135, 32'sd549, 32'sd1833,
32'sd513, 32'sd653, 32'sd1853, 32'sd1622, 32'sd917, 32'sd498,
32'sd1780, 32'sd1534, 32'sd645, 32'sd1743, 32'sd460, 32'sd1617,
32'sd822, 32'sd549, 32'sd236, 32'sd427, 32'sd310, 32'sd1715,
32'sd1491, 32'sd1033, 32'sd1044, 32'sd914, 32'sd739, 32'sd1644,
32'sd826, 32'sd1255, 32'sd1561, 32'sd1715, 32'sd591, 32'sd897,
32'sd340, 32'sd781, 32'sd618, 32'sd416, 32'sd671, 32'sd1248,
32'sd1066, 32'sd1605, 32'sd740, 32'sd1313, 32'sd1057, 32'sd450,
32'sd1103, 32'sd911, 32'sd1392, 32'sd233, 32'sd948, 32'sd278,
32'sd727, 32'sd783, 32'sd955, 32'sd1751, 32'sd322, 32'sd302,
32'sd830, 32'sd1989, 32'sd1115, 32'sd1812, 32'sd693, 32'sd1397,
32'sd157, 32'sd166, 32'sd1209, 32'sd1286, 32'sd372, 32'sd646,
32'sd298, 32'sd1049, 32'sd240, 32'sd1075, 32'sd1554, 32'sd771,
32'sd1315, 32'sd1139, 32'sd476, 32'sd1941, 32'sd531, 32'sd1267,
32'sd304, 32'sd1444, 32'sd1007, 32'sd877, 32'sd1689, 32'sd845,
32'sd212, 32'sd1401, 32'sd1452, 32'sd104, 32'sd986, 32'sd976,
32'sd1470, 32'sd1019, 32'sd1251, 32'sd208, 32'sd387, 32'sd1634,
32'sd747, 32'sd169, 32'sd958, 32'sd1762, 32'sd581, 32'sd1662,
32'sd1759, 32'sd1912, 32'sd1426, 32'sd516, 32'sd1816, 32'sd1152,
32'sd483, 32'sd1114, 32'sd1820, 32'sd1319, 32'sd1378, 32'sd1070,
32'sd750, 32'sd1557, 32'sd1879, 32'sd1792, 32'sd1438, 32'sd1409,
32'sd1619, 32'sd1392, 32'sd1168, 32'sd1627, 32'sd1845, 32'sd1923,
32'sd210, 32'sd1902, 32'sd1822, 32'sd517, 32'sd1149, 32'sd613,
32'sd1558, 32'sd1531, 32'sd1543, 32'sd699, 32'sd200, 32'sd1803,
32'sd1740, 32'sd1230, 32'sd1035, 32'sd1242, 32'sd1056, 32'sd952,
32'sd837, 32'sd1461, 32'sd512, 32'sd1934, 32'sd1740, 32'sd1583,
32'sd1884, 32'sd356, 32'sd1720, 32'sd956, 32'sd619, 32'sd554,
32'sd1164, 32'sd766, 32'sd1598, 32'sd1802, 32'sd560, 32'sd899,
32'sd635, 32'sd1915, 32'sd715, 32'sd1776, 32'sd533, 32'sd1768,
32'sd930, 32'sd232, 32'sd701, 32'sd910, 32'sd1270, 32'sd1365,
32'sd1233, 32'sd1365, 32'sd1950, 32'sd1083, 32'sd1001, 32'sd370,
32'sd914, 32'sd399, 32'sd1296, 32'sd1373, 32'sd1201, 32'sd289,
32'sd1211, 32'sd1407, 32'sd434, 32'sd1383, 32'sd291, 32'sd148,
32'sd210, 32'sd911, 32'sd147, 32'sd1436, 32'sd1527, 32'sd1898,
32'sd1300, 32'sd511, 32'sd126, 32'sd400, 32'sd158, 32'sd139,
32'sd925, 32'sd202, 32'sd549, 32'sd642, 32'sd234, 32'sd356,
32'sd1686, 32'sd1837, 32'sd1931, 32'sd171, 32'sd611, 32'sd1846,
32'sd633, 32'sd330, 32'sd1845, 32'sd1841, 32'sd1818, 32'sd122,
32'sd1508, 32'sd1550, 32'sd742, 32'sd698, 32'sd616, 32'sd1455,
32'sd607, 32'sd118, 32'sd1508, 32'sd852, 32'sd401, 32'sd1453,
32'sd742, 32'sd1289, 32'sd117, 32'sd1034, 32'sd939, 32'sd448,
32'sd1568, 32'sd100, 32'sd302, 32'sd864, 32'sd353, 32'sd1244,
32'sd1659, 32'sd669, 32'sd476, 32'sd210, 32'sd829, 32'sd1558,
32'sd550, 32'sd281, 32'sd1466, 32'sd1604, 32'sd439, 32'sd1447,
32'sd1408, 32'sd165, 32'sd526, 32'sd1928, 32'sd675, 32'sd187,
32'sd1466, 32'sd441, 32'sd734, 32'sd884, 32'sd685, 32'sd1982,
32'sd245, 32'sd1456, 32'sd1155, 32'sd1339, 32'sd1225, 32'sd1693,
32'sd794, 32'sd918, 32'sd679, 32'sd1898, 32'sd1002, 32'sd1438,
32'sd535, 32'sd756, 32'sd257, 32'sd242, 32'sd1072, 32'sd1460,
32'sd842, 32'sd617, 32'sd307, 32'sd1725, 32'sd1081, 32'sd1014,
32'sd311, 32'sd1454, 32'sd1543, 32'sd1431, 32'sd1839, 32'sd1590,
32'sd782, 32'sd537, 32'sd429, 32'sd455, 32'sd1414, 32'sd703,
32'sd1717, 32'sd1968, 32'sd787, 32'sd144, 32'sd773, 32'sd1925,
32'sd607, 32'sd159, 32'sd311, 32'sd1070, 32'sd1793, 32'sd1765,
32'sd731, 32'sd1645, 32'sd434, 32'sd961, 32'sd1668, 32'sd1263,
32'sd747, 32'sd683, 32'sd1599, 32'sd1918, 32'sd1981, 32'sd332,
32'sd675, 32'sd321, 32'sd1635, 32'sd831, 32'sd1124, 32'sd222,
32'sd1299, 32'sd1186, 32'sd1616, 32'sd562, 32'sd963, 32'sd1437,
32'sd504, 32'sd346, 32'sd1959, 32'sd1382, 32'sd331, 32'sd914,
32'sd575, 32'sd447, 32'sd1994, 32'sd1510, 32'sd1901, 32'sd1033,
32'sd639, 32'sd162, 32'sd346, 32'sd556, 32'sd1391, 32'sd758,
32'sd1481, 32'sd962, 32'sd1281, 32'sd1334, 32'sd1327, 32'sd1966,
32'sd1013, 32'sd1497, 32'sd934, 32'sd767, 32'sd1391, 32'sd1285,
32'sd1658, 32'sd774, 32'sd1239, 32'sd604, 32'sd1454, 32'sd172,
32'sd395, 32'sd965, 32'sd1458, 32'sd666, 32'sd142, 32'sd1423,
32'sd1998, 32'sd1787, 32'sd570, 32'sd1110, 32'sd1157, 32'sd940,
32'sd670, 32'sd422, 32'sd1733, 32'sd583, 32'sd518, 32'sd1516,
32'sd123, 32'sd1039, 32'sd1322, 32'sd1098, 32'sd965, 32'sd1419,
32'sd1153, 32'sd1442, 32'sd595, 32'sd1328, 32'sd642, 32'sd504,
32'sd1145, 32'sd948, 32'sd985, 32'sd1510, 32'sd1769, 32'sd187,
32'sd1932, 32'sd103, 32'sd1163, 32'sd386, 32'sd245, 32'sd1082,
32'sd882, 32'sd735, 32'sd947, 32'sd575, 32'sd916, 32'sd1449,
32'sd397, 32'sd1352, 32'sd909, 32'sd716, 32'sd1024, 32'sd1835,
32'sd635, 32'sd1405, 32'sd742, 32'sd1905, 32'sd859, 32'sd621,
32'sd1047, 32'sd1367, 32'sd741, 32'sd1995, 32'sd917, 32'sd1372,
32'sd1470, 32'sd1042, 32'sd1025, 32'sd586, 32'sd163, 32'sd563,
32'sd325, 32'sd1554, 32'sd1769, 32'sd1268, 32'sd768, 32'sd895,
32'sd581, 32'sd1671, 32'sd1227, 32'sd1445, 32'sd781, 32'sd218,
32'sd1444, 32'sd1836, 32'sd1540, 32'sd359, 32'sd709, 32'sd1294,
32'sd600, 32'sd592, 32'sd1369, 32'sd550, 32'sd307, 32'sd1819,
32'sd1300, 32'sd1055, 32'sd686, 32'sd768, 32'sd108, 32'sd1621,
32'sd1564, 32'sd631, 32'sd305, 32'sd1272, 32'sd139, 32'sd942,
32'sd890, 32'sd1367, 32'sd299, 32'sd1747, 32'sd1210, 32'sd1349,
32'sd350, 32'sd1918, 32'sd559, 32'sd1484, 32'sd1010, 32'sd628,
32'sd1697, 32'sd1589, 32'sd727, 32'sd789, 32'sd1805, 32'sd1659,
32'sd1298, 32'sd389, 32'sd910, 32'sd1105, 32'sd278, 32'sd1251,
32'sd1878, 32'sd1910, 32'sd597, 32'sd1664, 32'sd806, 32'sd1279,
32'sd1073, 32'sd1901, 32'sd576, 32'sd789, 32'sd1977, 32'sd1497,
32'sd169, 32'sd1972, 32'sd1719, 32'sd503, 32'sd1845, 32'sd1393,
32'sd413, 32'sd1787, 32'sd1631, 32'sd286, 32'sd250, 32'sd1785,
32'sd914, 32'sd808, 32'sd1738, 32'sd1635, 32'sd631, 32'sd142,
32'sd1770, 32'sd1047, 32'sd1067, 32'sd457, 32'sd1193, 32'sd1362,
32'sd507, 32'sd1548, 32'sd1978, 32'sd1243, 32'sd1599, 32'sd411,
32'sd305, 32'sd1708, 32'sd1572, 32'sd1030, 32'sd1867, 32'sd1114,
32'sd1125, 32'sd1768, 32'sd1640, 32'sd1193, 32'sd1312, 32'sd652,
32'sd833, 32'sd1640, 32'sd586, 32'sd1179, 32'sd1345, 32'sd354,
32'sd124, 32'sd1194, 32'sd1571, 32'sd324, 32'sd548, 32'sd722,
32'sd1224, 32'sd374, 32'sd1261, 32'sd1817, 32'sd554, 32'sd776,
32'sd1308, 32'sd614, 32'sd529, 32'sd1487, 32'sd982, 32'sd1845,
32'sd779, 32'sd1850, 32'sd1743, 32'sd924, 32'sd601, 32'sd1335,
32'sd743, 32'sd1394, 32'sd1675, 32'sd634, 32'sd1483, 32'sd736,
32'sd176, 32'sd1101, 32'sd1565, 32'sd623, 32'sd1198, 32'sd703,
32'sd1722, 32'sd918, 32'sd1234, 32'sd1354, 32'sd1414, 32'sd1265,
32'sd1362, 32'sd547, 32'sd568, 32'sd844, 32'sd1400, 32'sd199,
32'sd243, 32'sd302, 32'sd319, 32'sd1003, 32'sd733, 32'sd561,
32'sd284, 32'sd1678, 32'sd316, 32'sd814, 32'sd800, 32'sd601,
32'sd1694, 32'sd126, 32'sd1974, 32'sd331, 32'sd336, 32'sd978,
32'sd808, 32'sd178, 32'sd971, 32'sd419, 32'sd222, 32'sd991,
32'sd1854, 32'sd1745, 32'sd1502, 32'sd1305, 32'sd113, 32'sd1737,
32'sd912, 32'sd1463, 32'sd1950, 32'sd797, 32'sd1022, 32'sd1805,
32'sd1584, 32'sd700, 32'sd1910, 32'sd675, 32'sd1629, 32'sd1423,
32'sd289, 32'sd1451, 32'sd1915, 32'sd1986, 32'sd774, 32'sd1606,
32'sd1195, 32'sd152, 32'sd255, 32'sd203, 32'sd1830, 32'sd1937,
32'sd301, 32'sd785, 32'sd1160, 32'sd1491, 32'sd1431, 32'sd787,
32'sd1617, 32'sd988, 32'sd1619, 32'sd1745, 32'sd1640, 32'sd951,
32'sd1543, 32'sd1031, 32'sd380, 32'sd1042, 32'sd750, 32'sd445,
32'sd228, 32'sd312, 32'sd1513, 32'sd1045, 32'sd1776, 32'sd1403,
32'sd229, 32'sd442, 32'sd1565, 32'sd1038, 32'sd248, 32'sd1563,
32'sd1236, 32'sd1675, 32'sd682, 32'sd1958, 32'sd1915, 32'sd502,
32'sd446, 32'sd750, 32'sd143, 32'sd482, 32'sd1472, 32'sd1623,
32'sd947, 32'sd1644, 32'sd449, 32'sd1565, 32'sd437, 32'sd693,
32'sd176, 32'sd1295, 32'sd1962, 32'sd836, 32'sd842, 32'sd1038,
32'sd1328, 32'sd957, 32'sd673, 32'sd1225, 32'sd1144, 32'sd1523,
32'sd633, 32'sd1271, 32'sd1380, 32'sd911, 32'sd397, 32'sd1942,
32'sd1474, 32'sd1761, 32'sd1428, 32'sd891, 32'sd359, 32'sd182,
32'sd709, 32'sd513, 32'sd1782, 32'sd1876, 32'sd806, 32'sd1131,
32'sd1768, 32'sd1700, 32'sd543, 32'sd116, 32'sd1128, 32'sd1076,
32'sd656, 32'sd202, 32'sd1166, 32'sd596, 32'sd1960, 32'sd1058,
32'sd1020, 32'sd1563, 32'sd898, 32'sd1434, 32'sd1675, 32'sd1237,
32'sd1570, 32'sd344, 32'sd788, 32'sd1780, 32'sd1317, 32'sd944,
32'sd996, 32'sd1169, 32'sd1198, 32'sd391, 32'sd208, 32'sd1571,
32'sd1600, 32'sd648, 32'sd624, 32'sd286, 32'sd1400, 32'sd1404,
32'sd558, 32'sd306, 32'sd681, 32'sd1153, 32'sd1853, 32'sd326,
32'sd581, 32'sd1476, 32'sd496, 32'sd1179, 32'sd858, 32'sd206,
32'sd1108, 32'sd1116, 32'sd836, 32'sd194, 32'sd129, 32'sd1744,
32'sd1859, 32'sd1152, 32'sd1086, 32'sd1557, 32'sd426, 32'sd385,
32'sd397, 32'sd1280, 32'sd1637, 32'sd1845, 32'sd1418, 32'sd1349,
32'sd378, 32'sd1168, 32'sd265, 32'sd217, 32'sd1224, 32'sd1153,
32'sd1444, 32'sd1423, 32'sd635, 32'sd1551, 32'sd825, 32'sd336,
32'sd1381, 32'sd1239, 32'sd1292, 32'sd1866, 32'sd1650, 32'sd1160,
32'sd1944, 32'sd1129, 32'sd1860, 32'sd1603, 32'sd1742, 32'sd1280,
32'sd233, 32'sd740, 32'sd1941, 32'sd312, 32'sd274, 32'sd898,
32'sd968, 32'sd1827, 32'sd139, 32'sd1415, 32'sd813, 32'sd1854,
32'sd277, 32'sd1532, 32'sd1017, 32'sd512, 32'sd1597, 32'sd419,
32'sd568, 32'sd163, 32'sd987, 32'sd1540, 32'sd1083, 32'sd1430,
32'sd1790, 32'sd1000, 32'sd1771, 32'sd692, 32'sd651, 32'sd1946,
32'sd552, 32'sd1947, 32'sd1060, 32'sd1783, 32'sd1490, 32'sd1045,
32'sd622, 32'sd525, 32'sd689, 32'sd997, 32'sd1966, 32'sd727,
32'sd1109, 32'sd436, 32'sd914, 32'sd1217, 32'sd1846, 32'sd711,
32'sd918, 32'sd1649, 32'sd736, 32'sd510, 32'sd103, 32'sd208,
32'sd1678, 32'sd261, 32'sd1866, 32'sd876, 32'sd285, 32'sd1229,
32'sd1896, 32'sd1956, 32'sd1394, 32'sd1786, 32'sd1883, 32'sd691,
32'sd1322, 32'sd1246, 32'sd650, 32'sd919, 32'sd925, 32'sd1582,
32'sd1519, 32'sd1021, 32'sd1618, 32'sd1777, 32'sd1201, 32'sd1515,
32'sd1136, 32'sd917, 32'sd1369, 32'sd1878, 32'sd541, 32'sd1271,
32'sd990, 32'sd1138, 32'sd1913, 32'sd1253, 32'sd1440, 32'sd794,
32'sd1315, 32'sd472, 32'sd1616, 32'sd655, 32'sd1534, 32'sd158,
32'sd429, 32'sd930, 32'sd1294, 32'sd1548, 32'sd1860, 32'sd136,
32'sd1337, 32'sd1055, 32'sd997, 32'sd988, 32'sd797, 32'sd604,
32'sd765, 32'sd439, 32'sd1360, 32'sd314, 32'sd350, 32'sd1560,
32'sd439, 32'sd829, 32'sd546, 32'sd1471, 32'sd1481, 32'sd1706,
32'sd202, 32'sd863, 32'sd934, 32'sd917, 32'sd436, 32'sd341,
32'sd333, 32'sd707, 32'sd696, 32'sd1981, 32'sd1374, 32'sd1373,
32'sd122, 32'sd1784, 32'sd1969, 32'sd302, 32'sd266, 32'sd616,
32'sd1737, 32'sd850, 32'sd808, 32'sd1554, 32'sd713, 32'sd1919,
32'sd988, 32'sd1078, 32'sd1467, 32'sd1798, 32'sd928, 32'sd1665,
32'sd1441, 32'sd1692, 32'sd428, 32'sd1275, 32'sd158, 32'sd1674,
32'sd149, 32'sd1721, 32'sd1430, 32'sd1791, 32'sd493, 32'sd1346,
32'sd382, 32'sd1225, 32'sd976, 32'sd1299, 32'sd1293, 32'sd1562,
32'sd1965, 32'sd1378, 32'sd626, 32'sd1607, 32'sd304, 32'sd1770,
32'sd1608, 32'sd743, 32'sd981, 32'sd1367, 32'sd599, 32'sd1761,
32'sd1330, 32'sd447, 32'sd450, 32'sd112, 32'sd1572, 32'sd287,
32'sd746, 32'sd1989, 32'sd1993, 32'sd1208, 32'sd667, 32'sd881,
32'sd707, 32'sd1838, 32'sd887, 32'sd123, 32'sd648, 32'sd1852,
32'sd1606, 32'sd1425, 32'sd355, 32'sd1787, 32'sd1045, 32'sd307,
32'sd1608, 32'sd1629, 32'sd1853, 32'sd1044, 32'sd1469, 32'sd761,
32'sd909, 32'sd1490, 32'sd761, 32'sd839, 32'sd913, 32'sd1401,
32'sd1447, 32'sd471, 32'sd443, 32'sd1392, 32'sd1352, 32'sd1853,
32'sd1535, 32'sd1291, 32'sd161, 32'sd1862, 32'sd744, 32'sd1932,
32'sd920, 32'sd1368, 32'sd1978, 32'sd519, 32'sd814, 32'sd1425,
32'sd419, 32'sd936, 32'sd1291, 32'sd1546, 32'sd1606, 32'sd209,
32'sd1157, 32'sd1517, 32'sd252, 32'sd344, 32'sd790, 32'sd975,
32'sd1808, 32'sd1040, 32'sd1800, 32'sd360, 32'sd712, 32'sd398,
32'sd1403, 32'sd1504, 32'sd1227, 32'sd398, 32'sd816, 32'sd1855,
32'sd919, 32'sd1161, 32'sd556, 32'sd1789, 32'sd710, 32'sd1067,
32'sd1530, 32'sd497, 32'sd1235, 32'sd1974, 32'sd1706, 32'sd382,
32'sd757, 32'sd666, 32'sd869, 32'sd1903, 32'sd526, 32'sd1645,
32'sd1048, 32'sd1856, 32'sd252, 32'sd1534, 32'sd1084, 32'sd1055,
32'sd128, 32'sd278, 32'sd1784, 32'sd1720, 32'sd476, 32'sd1064,
32'sd1728, 32'sd1949, 32'sd1790, 32'sd1028, 32'sd1378, 32'sd324,
32'sd1316, 32'sd498, 32'sd1255, 32'sd1267, 32'sd397, 32'sd617,
32'sd1674, 32'sd324, 32'sd1305, 32'sd679, 32'sd886, 32'sd1427,
32'sd134, 32'sd263, 32'sd489, 32'sd1814, 32'sd1557, 32'sd1198,
32'sd1814, 32'sd819, 32'sd974, 32'sd1701, 32'sd474, 32'sd1241,
32'sd661, 32'sd485, 32'sd1565, 32'sd1538, 32'sd1168, 32'sd557,
32'sd1364, 32'sd1611, 32'sd454, 32'sd749, 32'sd798, 32'sd111,
32'sd1642, 32'sd726, 32'sd466, 32'sd1086, 32'sd1065, 32'sd1674,
32'sd1307, 32'sd817, 32'sd1768, 32'sd266, 32'sd1562, 32'sd1626,
32'sd942, 32'sd1517, 32'sd1613, 32'sd1656, 32'sd224, 32'sd1451,
32'sd1138, 32'sd1539, 32'sd155, 32'sd1913, 32'sd245, 32'sd985,
32'sd1226, 32'sd1828, 32'sd986, 32'sd197, 32'sd1143, 32'sd189,
32'sd1986, 32'sd1163, 32'sd532, 32'sd1419, 32'sd208, 32'sd1573,
32'sd222, 32'sd1151, 32'sd920, 32'sd1083, 32'sd992, 32'sd929,
32'sd1008, 32'sd1720, 32'sd775, 32'sd1217, 32'sd514, 32'sd754,
32'sd886, 32'sd1979, 32'sd1175, 32'sd1256, 32'sd1688, 32'sd788,
32'sd234, 32'sd1876, 32'sd500, 32'sd1648, 32'sd714, 32'sd1775,
32'sd328, 32'sd1062, 32'sd682, 32'sd219, 32'sd698, 32'sd930,
32'sd585, 32'sd1910, 32'sd583, 32'sd1979, 32'sd1407, 32'sd1630,
32'sd1537, 32'sd1190, 32'sd355, 32'sd388, 32'sd896, 32'sd1737,
32'sd1944, 32'sd245, 32'sd1317, 32'sd1650, 32'sd1181, 32'sd367,
32'sd167, 32'sd1796, 32'sd1773, 32'sd178, 32'sd568, 32'sd694,
32'sd1208, 32'sd1657, 32'sd346, 32'sd1525, 32'sd1055, 32'sd245,
32'sd878, 32'sd983, 32'sd1470, 32'sd1151, 32'sd1929, 32'sd1399,
32'sd890, 32'sd407, 32'sd945, 32'sd1664, 32'sd283, 32'sd1780,
32'sd205, 32'sd1491, 32'sd602, 32'sd128, 32'sd255, 32'sd1392,
32'sd1832, 32'sd520, 32'sd236, 32'sd1213, 32'sd846, 32'sd210,
32'sd647, 32'sd565, 32'sd1084, 32'sd119, 32'sd1581, 32'sd1471,
32'sd1561, 32'sd832, 32'sd1012, 32'sd429, 32'sd1060, 32'sd1436,
32'sd355, 32'sd1948, 32'sd1064, 32'sd481, 32'sd1426, 32'sd1998,
32'sd1636, 32'sd1604, 32'sd1885, 32'sd577, 32'sd1739, 32'sd837,
32'sd1004, 32'sd887, 32'sd1457, 32'sd1501, 32'sd515, 32'sd1510,
32'sd1716, 32'sd1151, 32'sd1092, 32'sd1728, 32'sd1524, 32'sd884,
32'sd1543, 32'sd619, 32'sd1127, 32'sd1452, 32'sd1771, 32'sd1033,
32'sd1731, 32'sd1698, 32'sd636, 32'sd1242, 32'sd1713, 32'sd1994,
32'sd1542, 32'sd1035, 32'sd1156, 32'sd397, 32'sd578, 32'sd564,
32'sd983, 32'sd1524, 32'sd1798, 32'sd1732, 32'sd1184, 32'sd536,
32'sd1098, 32'sd1406, 32'sd397, 32'sd563, 32'sd767, 32'sd291,
32'sd927, 32'sd1387, 32'sd186, 32'sd136, 32'sd1654, 32'sd883,
32'sd1489, 32'sd709, 32'sd838, 32'sd1583, 32'sd1741, 32'sd1942,
32'sd589, 32'sd1256, 32'sd398, 32'sd1670, 32'sd525, 32'sd486,
32'sd480, 32'sd732, 32'sd537, 32'sd833, 32'sd254, 32'sd1528,
32'sd487, 32'sd1162, 32'sd932, 32'sd1297, 32'sd1402, 32'sd1386,
32'sd1349, 32'sd1239, 32'sd1120, 32'sd726, 32'sd1288, 32'sd1479,
32'sd721, 32'sd543, 32'sd1724, 32'sd937, 32'sd178, 32'sd1015,
32'sd1116, 32'sd1456, 32'sd1747, 32'sd1198, 32'sd530, 32'sd1989,
32'sd687, 32'sd1392, 32'sd949, 32'sd176, 32'sd1079, 32'sd700,
32'sd296, 32'sd292, 32'sd1451, 32'sd1382, 32'sd360, 32'sd1061,
32'sd872, 32'sd886, 32'sd1305, 32'sd643, 32'sd1859, 32'sd1545,
32'sd625, 32'sd478, 32'sd677, 32'sd1402, 32'sd1701, 32'sd326,
32'sd431, 32'sd472, 32'sd633, 32'sd389, 32'sd584, 32'sd1982,
32'sd1475, 32'sd214, 32'sd1124, 32'sd894, 32'sd1522, 32'sd242,
32'sd1779, 32'sd1430, 32'sd1101, 32'sd172, 32'sd1007, 32'sd1378,
32'sd637, 32'sd1234, 32'sd185, 32'sd1380, 32'sd835, 32'sd753,
32'sd878, 32'sd1218, 32'sd1423, 32'sd333, 32'sd385, 32'sd1254,
32'sd451, 32'sd930, 32'sd113, 32'sd439, 32'sd1393, 32'sd1012,
32'sd1845, 32'sd610, 32'sd846, 32'sd1196, 32'sd287, 32'sd227,
32'sd863, 32'sd785, 32'sd1557, 32'sd482, 32'sd353, 32'sd974,
32'sd1544, 32'sd1559, 32'sd754, 32'sd1827, 32'sd289, 32'sd784,
32'sd357, 32'sd467, 32'sd1976, 32'sd1904, 32'sd1898, 32'sd833,
32'sd351, 32'sd1587, 32'sd1406, 32'sd1897, 32'sd1437, 32'sd522,
32'sd286, 32'sd1821, 32'sd1875, 32'sd1440, 32'sd1408, 32'sd1235,
32'sd729, 32'sd1981, 32'sd1880, 32'sd1218, 32'sd1503, 32'sd1384,
32'sd570, 32'sd1132, 32'sd943, 32'sd1938, 32'sd948, 32'sd473,
32'sd343, 32'sd783, 32'sd466, 32'sd269, 32'sd1493, 32'sd1236,
32'sd1928, 32'sd523, 32'sd1464, 32'sd340, 32'sd179, 32'sd478,
32'sd1667, 32'sd1020, 32'sd1678, 32'sd562, 32'sd1732, 32'sd223,
32'sd419, 32'sd741, 32'sd1439, 32'sd464, 32'sd1241, 32'sd1956,
32'sd480, 32'sd1982, 32'sd1072, 32'sd753, 32'sd152, 32'sd582,
32'sd539, 32'sd245, 32'sd1731, 32'sd495, 32'sd921, 32'sd240,
32'sd1020, 32'sd662, 32'sd253, 32'sd342, 32'sd586, 32'sd169,
32'sd625, 32'sd409, 32'sd773, 32'sd1944, 32'sd1852, 32'sd909,
32'sd704, 32'sd1885, 32'sd759, 32'sd1691, 32'sd1243, 32'sd914,
32'sd620, 32'sd1114, 32'sd1959, 32'sd119, 32'sd903, 32'sd1840,
32'sd1400, 32'sd777, 32'sd976, 32'sd911, 32'sd1769, 32'sd1650,
32'sd477, 32'sd1096, 32'sd202, 32'sd238, 32'sd934, 32'sd1686,
32'sd658, 32'sd1916, 32'sd1843, 32'sd543, 32'sd1768, 32'sd200,
32'sd1134, 32'sd183, 32'sd1873, 32'sd185, 32'sd1555, 32'sd1414,
32'sd725, 32'sd385, 32'sd1512, 32'sd495, 32'sd105, 32'sd1958,
32'sd1872, 32'sd392, 32'sd1979, 32'sd1001, 32'sd1069, 32'sd429,
32'sd1970, 32'sd1669, 32'sd1812, 32'sd1521, 32'sd707, 32'sd344,
32'sd1270, 32'sd541, 32'sd169, 32'sd504, 32'sd1483, 32'sd1289,
32'sd678, 32'sd1961, 32'sd905, 32'sd1121, 32'sd898, 32'sd1379,
32'sd303, 32'sd1813, 32'sd1579, 32'sd1702, 32'sd267, 32'sd778,
32'sd519, 32'sd920, 32'sd501, 32'sd1651, 32'sd1200, 32'sd847,
32'sd1047, 32'sd616, 32'sd517, 32'sd1246, 32'sd172, 32'sd1989,
32'sd1755, 32'sd133, 32'sd1455, 32'sd1315, 32'sd358, 32'sd1419,
32'sd1022, 32'sd1187, 32'sd986, 32'sd1236, 32'sd858, 32'sd994,
32'sd244, 32'sd1123, 32'sd299, 32'sd1429, 32'sd1855, 32'sd1237,
32'sd119, 32'sd1312, 32'sd280, 32'sd1617, 32'sd398, 32'sd1849,
32'sd1980, 32'sd279, 32'sd574, 32'sd1498, 32'sd243, 32'sd1813,
32'sd1938, 32'sd1876, 32'sd755, 32'sd1706, 32'sd557, 32'sd128,
32'sd1224, 32'sd475, 32'sd1151, 32'sd1922, 32'sd1506, 32'sd1694,
32'sd1152, 32'sd531, 32'sd379, 32'sd1219, 32'sd1782, 32'sd698,
32'sd717, 32'sd1148, 32'sd1730, 32'sd833, 32'sd720, 32'sd1777,
32'sd1618, 32'sd1884, 32'sd816, 32'sd276, 32'sd927, 32'sd827,
32'sd247, 32'sd885, 32'sd207, 32'sd899, 32'sd749, 32'sd1594,
32'sd911, 32'sd840, 32'sd1527, 32'sd1192, 32'sd145, 32'sd812,
32'sd347, 32'sd1672, 32'sd1201, 32'sd560, 32'sd245, 32'sd489,
32'sd392, 32'sd1645, 32'sd1377, 32'sd1571, 32'sd1744, 32'sd1434,
32'sd1904, 32'sd851, 32'sd349, 32'sd512, 32'sd1083, 32'sd1918,
32'sd1964, 32'sd1939, 32'sd304, 32'sd1294, 32'sd1449, 32'sd241,
32'sd1295, 32'sd1983, 32'sd501, 32'sd1054, 32'sd575, 32'sd1578,
32'sd262, 32'sd1854, 32'sd1912, 32'sd963, 32'sd1051, 32'sd930,
32'sd212, 32'sd393, 32'sd1716, 32'sd1942, 32'sd1841, 32'sd1510,
32'sd1211, 32'sd1873, 32'sd1990, 32'sd901, 32'sd335, 32'sd262,
32'sd1359, 32'sd1987, 32'sd1527, 32'sd660, 32'sd1795, 32'sd1369,
32'sd1582, 32'sd1427, 32'sd1655, 32'sd574, 32'sd943, 32'sd1235,
32'sd1083, 32'sd752, 32'sd1684, 32'sd808, 32'sd1972, 32'sd1800,
32'sd1364, 32'sd1798, 32'sd1249, 32'sd1613, 32'sd802, 32'sd1082,
32'sd857, 32'sd175, 32'sd115, 32'sd1887, 32'sd1726, 32'sd1449,
32'sd1218, 32'sd1234, 32'sd777, 32'sd903, 32'sd1995, 32'sd465,
32'sd159, 32'sd1655, 32'sd1361, 32'sd1051, 32'sd1185, 32'sd1007,
32'sd1578, 32'sd911, 32'sd1039, 32'sd1539, 32'sd1946, 32'sd1707,
32'sd1540, 32'sd718, 32'sd1460, 32'sd1761, 32'sd1347, 32'sd188,
32'sd937, 32'sd401, 32'sd971, 32'sd984, 32'sd513, 32'sd975,
32'sd471, 32'sd1030, 32'sd228, 32'sd458, 32'sd1977, 32'sd919,
32'sd1362, 32'sd1374, 32'sd1360, 32'sd994, 32'sd724, 32'sd377,
32'sd850, 32'sd1273, 32'sd684, 32'sd176, 32'sd684, 32'sd1422,
32'sd471, 32'sd1932, 32'sd1559, 32'sd1150, 32'sd193, 32'sd1792,
32'sd1093, 32'sd976, 32'sd899, 32'sd1608, 32'sd1885, 32'sd541,
32'sd556, 32'sd1578, 32'sd1235, 32'sd764, 32'sd1320, 32'sd705,
32'sd1751, 32'sd1712, 32'sd1492, 32'sd990, 32'sd376, 32'sd1447,
32'sd1824, 32'sd772, 32'sd674, 32'sd699, 32'sd1784, 32'sd358,
32'sd1439, 32'sd712, 32'sd1240, 32'sd901, 32'sd693, 32'sd1509,
32'sd1421, 32'sd1405, 32'sd1869, 32'sd1072, 32'sd1515, 32'sd1008,
32'sd645, 32'sd126, 32'sd1405, 32'sd500, 32'sd1277, 32'sd977,
32'sd542, 32'sd1753, 32'sd796, 32'sd839, 32'sd1565, 32'sd126,
32'sd1545, 32'sd371, 32'sd1187, 32'sd1397, 32'sd1691, 32'sd975,
32'sd1891, 32'sd1127, 32'sd442, 32'sd823, 32'sd110, 32'sd1572,
32'sd762, 32'sd750, 32'sd1839, 32'sd1386, 32'sd960, 32'sd1301,
32'sd631, 32'sd912, 32'sd1260, 32'sd307, 32'sd763, 32'sd417,
32'sd1461, 32'sd1280, 32'sd1217, 32'sd1596, 32'sd1621, 32'sd1238,
32'sd1769, 32'sd1418, 32'sd1818, 32'sd231, 32'sd1268, 32'sd452,
32'sd514, 32'sd255, 32'sd478, 32'sd127, 32'sd1545, 32'sd175,
32'sd1542, 32'sd1609, 32'sd1696, 32'sd436, 32'sd257, 32'sd133,
32'sd1975, 32'sd1541, 32'sd1135, 32'sd1282, 32'sd669, 32'sd475,
32'sd1574, 32'sd758, 32'sd1960, 32'sd1251, 32'sd1157, 32'sd619,
32'sd159, 32'sd1028, 32'sd156, 32'sd1412, 32'sd832, 32'sd1016,
32'sd1185, 32'sd704, 32'sd218, 32'sd913, 32'sd1173, 32'sd989,
32'sd506, 32'sd1160, 32'sd1675, 32'sd1144, 32'sd1765, 32'sd1752,
32'sd1340, 32'sd630, 32'sd202, 32'sd385, 32'sd301, 32'sd1689,
32'sd787, 32'sd1242, 32'sd128, 32'sd851, 32'sd574, 32'sd314,
32'sd543, 32'sd809, 32'sd1334, 32'sd875, 32'sd1460, 32'sd1087,
32'sd277, 32'sd1029, 32'sd765, 32'sd423, 32'sd171, 32'sd1712,
32'sd501, 32'sd337, 32'sd727, 32'sd1304, 32'sd1798, 32'sd819,
32'sd1642, 32'sd1829, 32'sd1029, 32'sd1397, 32'sd1308, 32'sd1072,
32'sd1380, 32'sd519, 32'sd714, 32'sd1287, 32'sd1661, 32'sd226,
32'sd564, 32'sd774, 32'sd1198, 32'sd412, 32'sd182, 32'sd1477,
32'sd1361, 32'sd654, 32'sd1089, 32'sd958, 32'sd189, 32'sd1566,
32'sd1060, 32'sd1112, 32'sd371, 32'sd1389, 32'sd807, 32'sd1024,
32'sd947, 32'sd380, 32'sd1186, 32'sd467, 32'sd1748, 32'sd1364,
32'sd1333, 32'sd1749, 32'sd1996, 32'sd1441, 32'sd377, 32'sd717,
32'sd1887, 32'sd1172, 32'sd1600, 32'sd1810, 32'sd1626, 32'sd362,
32'sd1571, 32'sd607, 32'sd1271, 32'sd1565, 32'sd851, 32'sd472,
32'sd1079, 32'sd1808, 32'sd842, 32'sd1208, 32'sd422, 32'sd1340,
32'sd437, 32'sd906, 32'sd1996, 32'sd188, 32'sd126, 32'sd706,
32'sd1147, 32'sd1892, 32'sd112, 32'sd606, 32'sd1885, 32'sd1767,
32'sd1155, 32'sd147, 32'sd420, 32'sd530, 32'sd1095, 32'sd1700,
32'sd880, 32'sd1174, 32'sd1612, 32'sd1824, 32'sd1682, 32'sd1862,
32'sd1013, 32'sd615, 32'sd1865, 32'sd1930, 32'sd1849, 32'sd1247,
32'sd1663, 32'sd1634, 32'sd1755, 32'sd1238, 32'sd1225, 32'sd1751,
32'sd180, 32'sd1827, 32'sd715, 32'sd660, 32'sd908, 32'sd498,
32'sd531, 32'sd1984, 32'sd1397, 32'sd1799, 32'sd1819, 32'sd1971,
32'sd281, 32'sd875, 32'sd1814, 32'sd1206, 32'sd145, 32'sd249,
32'sd1844, 32'sd786, 32'sd681, 32'sd209, 32'sd678, 32'sd1785,
32'sd1772, 32'sd1083, 32'sd972, 32'sd874, 32'sd1920, 32'sd1170,
32'sd170, 32'sd727, 32'sd1815, 32'sd1953, 32'sd1507, 32'sd683,
32'sd684, 32'sd1671, 32'sd1255, 32'sd1432, 32'sd935, 32'sd871,
32'sd1437, 32'sd286, 32'sd984, 32'sd1469, 32'sd142, 32'sd905,
32'sd642, 32'sd1686, 32'sd1834, 32'sd887, 32'sd1063, 32'sd1968,
32'sd1020, 32'sd1202, 32'sd209, 32'sd1608, 32'sd1591, 32'sd483,
32'sd543, 32'sd1226, 32'sd1373, 32'sd1187, 32'sd891, 32'sd1842,
32'sd209, 32'sd203, 32'sd1926, 32'sd467, 32'sd1336, 32'sd480,
32'sd1429, 32'sd1124, 32'sd1064, 32'sd1594, 32'sd1773, 32'sd1359,
32'sd1636, 32'sd739, 32'sd814, 32'sd1398, 32'sd804, 32'sd383,
32'sd215, 32'sd1716, 32'sd1173, 32'sd694, 32'sd1511, 32'sd944,
32'sd886, 32'sd1565, 32'sd1410, 32'sd132, 32'sd1838, 32'sd1926,
32'sd1006, 32'sd425, 32'sd1663, 32'sd296, 32'sd1372, 32'sd1455,
32'sd235, 32'sd151, 32'sd1701, 32'sd1392, 32'sd1591, 32'sd1076,
32'sd940, 32'sd1473, 32'sd1236, 32'sd135, 32'sd347, 32'sd1756,
32'sd1699, 32'sd1115, 32'sd750, 32'sd480, 32'sd1706, 32'sd1379,
32'sd1203, 32'sd492, 32'sd1335, 32'sd1213, 32'sd1431, 32'sd1665,
32'sd1777, 32'sd816, 32'sd1931, 32'sd1938, 32'sd1431, 32'sd578,
32'sd1863, 32'sd1231, 32'sd439, 32'sd1394, 32'sd1084, 32'sd1146,
32'sd423, 32'sd1664, 32'sd1431, 32'sd1407, 32'sd1485, 32'sd1007,
32'sd1003, 32'sd345, 32'sd1442, 32'sd1330, 32'sd1610, 32'sd617,
32'sd616, 32'sd1078, 32'sd842, 32'sd1924, 32'sd795, 32'sd1574,
32'sd729, 32'sd1711, 32'sd1374, 32'sd858, 32'sd140, 32'sd1531,
32'sd554, 32'sd398, 32'sd498, 32'sd868, 32'sd804, 32'sd455,
32'sd352, 32'sd714, 32'sd1268, 32'sd1777, 32'sd523, 32'sd1085,
32'sd1409, 32'sd1979, 32'sd993, 32'sd1562, 32'sd944, 32'sd1746,
32'sd1302, 32'sd1316, 32'sd1651, 32'sd1230, 32'sd1144, 32'sd1028,
32'sd227, 32'sd1598, 32'sd1034, 32'sd1966, 32'sd615, 32'sd525,
32'sd390, 32'sd853, 32'sd1926, 32'sd862, 32'sd1595, 32'sd1056,
32'sd956, 32'sd500, 32'sd1883, 32'sd1921, 32'sd1091, 32'sd144,
32'sd509, 32'sd443, 32'sd1665, 32'sd783, 32'sd1598, 32'sd321,
32'sd625, 32'sd1528, 32'sd1102, 32'sd540, 32'sd886, 32'sd715,
32'sd686, 32'sd808, 32'sd1131, 32'sd1101, 32'sd230, 32'sd123,
32'sd1861, 32'sd1343, 32'sd332, 32'sd141, 32'sd1332, 32'sd828,
32'sd791, 32'sd160, 32'sd1712, 32'sd1340, 32'sd1072, 32'sd600,
32'sd354, 32'sd845, 32'sd1974, 32'sd946, 32'sd458, 32'sd107,
32'sd1493, 32'sd713, 32'sd179, 32'sd524, 32'sd804, 32'sd623,
32'sd867, 32'sd637, 32'sd242, 32'sd928, 32'sd996, 32'sd904,
32'sd930, 32'sd901, 32'sd343, 32'sd187, 32'sd1033, 32'sd1306,
32'sd816, 32'sd1077, 32'sd1373, 32'sd402, 32'sd854, 32'sd601,
32'sd814, 32'sd1680, 32'sd414, 32'sd1402, 32'sd1609, 32'sd1969,
32'sd1104, 32'sd734, 32'sd261, 32'sd915, 32'sd615, 32'sd1039,
32'sd999, 32'sd1337, 32'sd386, 32'sd558, 32'sd539, 32'sd200,
32'sd1543, 32'sd1804, 32'sd1661, 32'sd1960, 32'sd1898, 32'sd1031,
32'sd1371, 32'sd1563, 32'sd151, 32'sd1127, 32'sd1155, 32'sd1682,
32'sd1555, 32'sd1969, 32'sd106, 32'sd850, 32'sd1848, 32'sd1762,
32'sd1608, 32'sd1617, 32'sd1130, 32'sd1145, 32'sd1217, 32'sd106,
32'sd973, 32'sd1159, 32'sd1540, 32'sd589, 32'sd1782, 32'sd661,
32'sd1725, 32'sd337, 32'sd1905, 32'sd426, 32'sd247, 32'sd1273,
32'sd121, 32'sd432, 32'sd849, 32'sd634, 32'sd1976, 32'sd1942,
32'sd904, 32'sd1011, 32'sd1620, 32'sd934, 32'sd1383, 32'sd586,
32'sd1987, 32'sd1767, 32'sd1662, 32'sd774, 32'sd926, 32'sd875,
32'sd657, 32'sd1289, 32'sd495, 32'sd1442, 32'sd529, 32'sd893,
32'sd868, 32'sd1465, 32'sd1612, 32'sd1864, 32'sd1316, 32'sd1498,
32'sd1338, 32'sd1576, 32'sd1253, 32'sd477, 32'sd941, 32'sd1889,
32'sd1221, 32'sd1450, 32'sd577, 32'sd1610, 32'sd1576, 32'sd1381,
32'sd1349, 32'sd768, 32'sd232, 32'sd463, 32'sd1359, 32'sd1389,
32'sd1257, 32'sd157, 32'sd1559, 32'sd1078, 32'sd749, 32'sd1709,
32'sd477, 32'sd627, 32'sd1291, 32'sd312, 32'sd1820, 32'sd1844,
32'sd1713, 32'sd704, 32'sd1140, 32'sd502, 32'sd783, 32'sd379,
32'sd1492, 32'sd1704, 32'sd1444, 32'sd1524, 32'sd896, 32'sd409,
32'sd968, 32'sd1095, 32'sd958, 32'sd406, 32'sd847, 32'sd1703,
32'sd1037, 32'sd1652, 32'sd1773, 32'sd1253, 32'sd1829, 32'sd770,
32'sd1506, 32'sd742, 32'sd1489, 32'sd335, 32'sd1955, 32'sd1416,
32'sd1768, 32'sd1062, 32'sd1314, 32'sd463, 32'sd1944, 32'sd1270,
32'sd202, 32'sd815, 32'sd693, 32'sd1122, 32'sd647, 32'sd1805,
32'sd946, 32'sd1824, 32'sd600, 32'sd1841, 32'sd1263, 32'sd211,
32'sd1956, 32'sd563, 32'sd973, 32'sd318, 32'sd1193, 32'sd777,
32'sd596, 32'sd1108, 32'sd822, 32'sd1669, 32'sd1660, 32'sd441,
32'sd1901, 32'sd1630, 32'sd1752, 32'sd404, 32'sd1173, 32'sd1551,
32'sd236, 32'sd1499, 32'sd680, 32'sd1912, 32'sd1441, 32'sd1190,
32'sd480, 32'sd1834, 32'sd1669, 32'sd645, 32'sd641, 32'sd991,
32'sd1364, 32'sd369, 32'sd288, 32'sd1804, 32'sd552, 32'sd1006,
32'sd1483, 32'sd1661, 32'sd1121, 32'sd1817, 32'sd712, 32'sd736,
32'sd1484, 32'sd1489, 32'sd1322, 32'sd1098, 32'sd1978, 32'sd760,
32'sd1800, 32'sd793, 32'sd1465, 32'sd874, 32'sd1246, 32'sd1776,
32'sd1860, 32'sd1265, 32'sd528, 32'sd1835, 32'sd1300, 32'sd1657,
32'sd874, 32'sd587, 32'sd1234, 32'sd147, 32'sd679, 32'sd1491,
32'sd512, 32'sd973, 32'sd725, 32'sd1038, 32'sd1134, 32'sd885,
32'sd1531, 32'sd973, 32'sd516, 32'sd1196, 32'sd502, 32'sd1552,
32'sd1742, 32'sd403, 32'sd862, 32'sd457, 32'sd1472, 32'sd1444,
32'sd1721, 32'sd1525, 32'sd599, 32'sd1007, 32'sd223, 32'sd952,
32'sd1472, 32'sd766, 32'sd1081, 32'sd1032, 32'sd1180, 32'sd612,
32'sd1343, 32'sd1814, 32'sd1579, 32'sd1383, 32'sd1026, 32'sd769,
32'sd642, 32'sd830, 32'sd964, 32'sd1379, 32'sd885, 32'sd1080,
32'sd931, 32'sd838, 32'sd545, 32'sd1284, 32'sd226, 32'sd595,
32'sd185, 32'sd1063, 32'sd689, 32'sd193, 32'sd116, 32'sd1484,
32'sd170, 32'sd1586, 32'sd1595, 32'sd1644, 32'sd1959, 32'sd1566,
32'sd849, 32'sd1301, 32'sd729, 32'sd1037, 32'sd318, 32'sd1970,
32'sd672, 32'sd1858, 32'sd1547, 32'sd434, 32'sd1773, 32'sd890,
32'sd1993, 32'sd1539, 32'sd620, 32'sd1461, 32'sd1102, 32'sd1160,
32'sd1960, 32'sd848, 32'sd608, 32'sd857, 32'sd1708, 32'sd1803,
32'sd321, 32'sd1746, 32'sd1836, 32'sd784, 32'sd1604, 32'sd733,
32'sd1870, 32'sd1373, 32'sd170, 32'sd1109, 32'sd709, 32'sd354,
32'sd236, 32'sd305, 32'sd172, 32'sd1728, 32'sd238, 32'sd1630,
32'sd1454, 32'sd443, 32'sd992, 32'sd724, 32'sd431, 32'sd1825,
32'sd586, 32'sd1785, 32'sd939, 32'sd1076, 32'sd738, 32'sd1733,
32'sd1756, 32'sd1664, 32'sd163, 32'sd1625, 32'sd1615, 32'sd723,
32'sd709, 32'sd371, 32'sd627, 32'sd577, 32'sd1625, 32'sd1879,
32'sd1145, 32'sd685, 32'sd1530, 32'sd328, 32'sd442, 32'sd1966,
32'sd648, 32'sd1323, 32'sd1265, 32'sd366, 32'sd885, 32'sd951,
32'sd1560, 32'sd1895, 32'sd1559, 32'sd1356, 32'sd412, 32'sd1790,
32'sd209, 32'sd283, 32'sd924, 32'sd260, 32'sd896, 32'sd138,
32'sd1334, 32'sd1839, 32'sd1998, 32'sd1892, 32'sd716, 32'sd1373,
32'sd277, 32'sd1816, 32'sd1050, 32'sd273, 32'sd1155, 32'sd841,
32'sd464, 32'sd1527, 32'sd1653, 32'sd1817, 32'sd1261, 32'sd1654,
32'sd453, 32'sd1050, 32'sd1371, 32'sd1374, 32'sd1397, 32'sd1928,
32'sd1704, 32'sd128, 32'sd1662, 32'sd1173, 32'sd289, 32'sd132,
32'sd560, 32'sd188, 32'sd1159, 32'sd528, 32'sd581, 32'sd552,
32'sd609, 32'sd250, 32'sd1393, 32'sd218, 32'sd781, 32'sd1619,
32'sd886, 32'sd1055, 32'sd1556, 32'sd1857, 32'sd149, 32'sd787,
32'sd150, 32'sd625, 32'sd1800, 32'sd1747, 32'sd1759, 32'sd695,
32'sd297, 32'sd1978, 32'sd270, 32'sd927, 32'sd332, 32'sd1863,
32'sd1753, 32'sd1806, 32'sd292, 32'sd833, 32'sd1372, 32'sd184,
32'sd1101, 32'sd572, 32'sd379, 32'sd1189, 32'sd1068, 32'sd376,
32'sd119, 32'sd1355, 32'sd1084, 32'sd1751, 32'sd1383, 32'sd1837,
32'sd837, 32'sd364, 32'sd1756, 32'sd807, 32'sd600, 32'sd353,
32'sd997, 32'sd1650, 32'sd1031, 32'sd1699, 32'sd1289, 32'sd820,
32'sd558, 32'sd1163, 32'sd1226, 32'sd330, 32'sd1290, 32'sd622,
32'sd696, 32'sd1184, 32'sd681, 32'sd982, 32'sd1961, 32'sd369,
32'sd878, 32'sd150, 32'sd1568, 32'sd200, 32'sd1642, 32'sd1126,
32'sd541, 32'sd523, 32'sd287, 32'sd388, 32'sd1825, 32'sd940,
32'sd1035, 32'sd1278, 32'sd197, 32'sd700, 32'sd1256, 32'sd1996,
32'sd925, 32'sd774, 32'sd1276, 32'sd708, 32'sd398, 32'sd977,
32'sd615, 32'sd986, 32'sd1112, 32'sd626, 32'sd481, 32'sd646,
32'sd1033, 32'sd1083, 32'sd311, 32'sd607, 32'sd784, 32'sd1103,
32'sd1951, 32'sd1104, 32'sd820, 32'sd1151, 32'sd983, 32'sd973,
32'sd295, 32'sd253, 32'sd125, 32'sd854, 32'sd184, 32'sd115,
32'sd1791, 32'sd1013, 32'sd1638, 32'sd226, 32'sd449, 32'sd661,
32'sd510, 32'sd467, 32'sd1489, 32'sd1566, 32'sd745, 32'sd1685,
32'sd1265, 32'sd1870, 32'sd1982, 32'sd1990, 32'sd1570, 32'sd1892,
32'sd1721, 32'sd208, 32'sd785, 32'sd644, 32'sd1195, 32'sd1132,
32'sd740, 32'sd1454, 32'sd840, 32'sd1312, 32'sd132, 32'sd941,
32'sd1699, 32'sd1178, 32'sd581, 32'sd1155, 32'sd986, 32'sd100,
32'sd811, 32'sd454, 32'sd1090, 32'sd1599, 32'sd1543, 32'sd298,
32'sd439, 32'sd721, 32'sd1521, 32'sd950, 32'sd873, 32'sd555,
32'sd1846, 32'sd292, 32'sd1348, 32'sd1312, 32'sd1189, 32'sd1436,
32'sd1879, 32'sd332, 32'sd922, 32'sd336, 32'sd501, 32'sd890,
32'sd128, 32'sd223, 32'sd1968, 32'sd537, 32'sd1128, 32'sd456,
32'sd453, 32'sd1779, 32'sd1698, 32'sd573, 32'sd447, 32'sd1056,
32'sd1906, 32'sd1488, 32'sd400, 32'sd1198, 32'sd1214, 32'sd1668,
32'sd430, 32'sd1359, 32'sd980, 32'sd990, 32'sd1159, 32'sd1429,
32'sd1175, 32'sd1743, 32'sd1684, 32'sd570, 32'sd1817, 32'sd109,
32'sd1661, 32'sd1723, 32'sd880, 32'sd1891, 32'sd709, 32'sd1447,
32'sd1260, 32'sd696, 32'sd1016, 32'sd883, 32'sd1288, 32'sd761,
32'sd473, 32'sd1268, 32'sd861, 32'sd1951, 32'sd1593, 32'sd475,
32'sd1501, 32'sd449, 32'sd1382, 32'sd718, 32'sd209, 32'sd385,
32'sd463, 32'sd929, 32'sd1680, 32'sd1009, 32'sd1944, 32'sd432,
32'sd1661, 32'sd253, 32'sd1423, 32'sd959, 32'sd671, 32'sd357,
32'sd380, 32'sd433, 32'sd1157, 32'sd728, 32'sd1287, 32'sd1271,
32'sd1911, 32'sd718, 32'sd148, 32'sd1185, 32'sd855, 32'sd305,
32'sd601, 32'sd332, 32'sd1573, 32'sd1201, 32'sd1220, 32'sd254,
32'sd1363, 32'sd692, 32'sd597, 32'sd368, 32'sd433, 32'sd1283,
32'sd717, 32'sd1152, 32'sd669, 32'sd1659, 32'sd405, 32'sd608,
32'sd1336, 32'sd1683, 32'sd1747, 32'sd1844, 32'sd139, 32'sd1722,
32'sd1024, 32'sd1169, 32'sd684, 32'sd1222, 32'sd1559, 32'sd1751,
32'sd983, 32'sd696, 32'sd1731, 32'sd885, 32'sd1449, 32'sd1511,
32'sd1717, 32'sd1555, 32'sd1500, 32'sd262, 32'sd906, 32'sd1759,
32'sd801, 32'sd1977, 32'sd458, 32'sd621, 32'sd1493, 32'sd1227,
32'sd1370, 32'sd365, 32'sd408, 32'sd510, 32'sd1897, 32'sd391,
32'sd1685, 32'sd895, 32'sd1599, 32'sd1238, 32'sd1277, 32'sd1392,
32'sd1804, 32'sd412, 32'sd1288, 32'sd186, 32'sd1844, 32'sd1889,
32'sd1790, 32'sd1564, 32'sd1852, 32'sd415, 32'sd887, 32'sd193,
32'sd1791, 32'sd592, 32'sd725, 32'sd194, 32'sd1254, 32'sd388,
32'sd780, 32'sd1196, 32'sd1606, 32'sd108, 32'sd1070, 32'sd931,
32'sd406, 32'sd807, 32'sd658, 32'sd1365, 32'sd101, 32'sd916,
32'sd1629, 32'sd819, 32'sd1595, 32'sd1663, 32'sd577, 32'sd1360,
32'sd101, 32'sd529, 32'sd449, 32'sd185, 32'sd1235, 32'sd420,
32'sd1713, 32'sd1084, 32'sd1518, 32'sd571, 32'sd859, 32'sd707,
32'sd1531, 32'sd1039, 32'sd173, 32'sd863, 32'sd736, 32'sd982,
32'sd585, 32'sd304, 32'sd1863, 32'sd238, 32'sd304, 32'sd903,
32'sd110, 32'sd1933, 32'sd356, 32'sd529, 32'sd801, 32'sd1131,
32'sd1127, 32'sd1393, 32'sd1342, 32'sd832, 32'sd411, 32'sd1960,
32'sd1890, 32'sd730, 32'sd430, 32'sd1034, 32'sd182, 32'sd1294,
32'sd1409, 32'sd691, 32'sd109, 32'sd1035, 32'sd593, 32'sd1458,
32'sd1351, 32'sd1839, 32'sd840, 32'sd1467, 32'sd1963, 32'sd831,
32'sd995, 32'sd1125, 32'sd1694, 32'sd367, 32'sd555, 32'sd1115,
32'sd107, 32'sd474, 32'sd1535, 32'sd1566, 32'sd1274, 32'sd1342,
32'sd901, 32'sd1079, 32'sd990, 32'sd516, 32'sd132, 32'sd573,
32'sd1762, 32'sd1543, 32'sd749, 32'sd1225, 32'sd1420, 32'sd501,
32'sd265, 32'sd1892, 32'sd579, 32'sd1401, 32'sd1719, 32'sd1101,
32'sd1616, 32'sd1128, 32'sd562, 32'sd1106, 32'sd652, 32'sd161,
32'sd261, 32'sd600, 32'sd1953, 32'sd1167, 32'sd149, 32'sd1994,
32'sd1676, 32'sd236, 32'sd1837, 32'sd1161, 32'sd1350, 32'sd1430,
32'sd1245, 32'sd130, 32'sd253, 32'sd184, 32'sd531, 32'sd1806,
32'sd279, 32'sd1570, 32'sd1778, 32'sd1274, 32'sd1507, 32'sd181,
32'sd1741, 32'sd1341, 32'sd451, 32'sd1682, 32'sd838, 32'sd1479,
32'sd615, 32'sd438, 32'sd1658, 32'sd612, 32'sd1589, 32'sd103,
32'sd1217, 32'sd667, 32'sd639, 32'sd882, 32'sd480, 32'sd1207,
32'sd920, 32'sd1070, 32'sd1198, 32'sd1311, 32'sd947, 32'sd1020,
32'sd1851, 32'sd956, 32'sd369, 32'sd1825, 32'sd358, 32'sd879,
32'sd877, 32'sd641, 32'sd183, 32'sd311, 32'sd258, 32'sd1540,
32'sd672, 32'sd387, 32'sd1661, 32'sd1300, 32'sd1790, 32'sd870,
32'sd158, 32'sd1042, 32'sd636, 32'sd919, 32'sd857, 32'sd1846,
32'sd1317, 32'sd1684, 32'sd409, 32'sd1574, 32'sd400, 32'sd670,
32'sd1980, 32'sd1230, 32'sd463, 32'sd159, 32'sd1112, 32'sd483,
32'sd480, 32'sd345, 32'sd599, 32'sd1738, 32'sd624, 32'sd563,
32'sd1425, 32'sd1838, 32'sd954, 32'sd1874, 32'sd264, 32'sd259,
32'sd1542, 32'sd1416, 32'sd1929, 32'sd1653, 32'sd466, 32'sd906,
32'sd829, 32'sd814, 32'sd1214, 32'sd801, 32'sd1422, 32'sd1531,
32'sd804, 32'sd1954, 32'sd330, 32'sd305, 32'sd1366, 32'sd1089,
32'sd1531, 32'sd1423, 32'sd1267, 32'sd442, 32'sd1632, 32'sd1227,
32'sd1839, 32'sd661, 32'sd1414, 32'sd151, 32'sd152, 32'sd280,
32'sd903, 32'sd1993, 32'sd1174, 32'sd1955, 32'sd757, 32'sd1033,
32'sd1487, 32'sd971, 32'sd1389, 32'sd1896, 32'sd852, 32'sd1117,
32'sd1748, 32'sd402, 32'sd502, 32'sd986, 32'sd202, 32'sd1671,
32'sd789, 32'sd1932, 32'sd1340, 32'sd1161, 32'sd419, 32'sd1155,
32'sd1403, 32'sd1255, 32'sd1564, 32'sd905, 32'sd1517, 32'sd1698,
32'sd1025, 32'sd1888, 32'sd409, 32'sd1874, 32'sd1718, 32'sd1833,
32'sd264, 32'sd1952, 32'sd1900, 32'sd1730, 32'sd449, 32'sd680,
32'sd450, 32'sd1016, 32'sd1290, 32'sd1854, 32'sd216, 32'sd584,
32'sd719, 32'sd1235, 32'sd1754, 32'sd241, 32'sd1593, 32'sd547,
32'sd1886, 32'sd147, 32'sd921, 32'sd1448, 32'sd809, 32'sd1023,
32'sd758, 32'sd745, 32'sd1223, 32'sd822, 32'sd1936, 32'sd501,
32'sd1927, 32'sd1208, 32'sd1931, 32'sd1938, 32'sd278, 32'sd322,
32'sd625, 32'sd747, 32'sd1484, 32'sd1790, 32'sd656, 32'sd540,
32'sd747, 32'sd506, 32'sd1202, 32'sd1841, 32'sd185, 32'sd1538,
32'sd1385, 32'sd1519, 32'sd883, 32'sd1482, 32'sd310, 32'sd1877,
32'sd361, 32'sd612, 32'sd1533, 32'sd1232, 32'sd1959, 32'sd1568,
32'sd1328, 32'sd1144, 32'sd1090, 32'sd1769, 32'sd836, 32'sd806,
32'sd1177, 32'sd1850, 32'sd1519, 32'sd1528, 32'sd664, 32'sd128,
32'sd802, 32'sd470, 32'sd645, 32'sd1897, 32'sd1338, 32'sd527,
32'sd1625, 32'sd1908, 32'sd1236, 32'sd1380, 32'sd1067, 32'sd771,
32'sd1230, 32'sd1254, 32'sd1079, 32'sd1652, 32'sd1065, 32'sd739,
32'sd936, 32'sd1720, 32'sd1346, 32'sd417, 32'sd566, 32'sd1489,
32'sd772, 32'sd1577, 32'sd968, 32'sd1685, 32'sd1669, 32'sd1339,
32'sd737, 32'sd1099, 32'sd1298, 32'sd1409, 32'sd823, 32'sd1571,
32'sd1594, 32'sd957, 32'sd1376, 32'sd958, 32'sd1315, 32'sd711,
32'sd1086, 32'sd211, 32'sd1528, 32'sd1622, 32'sd1350, 32'sd1073,
32'sd1676, 32'sd1394, 32'sd871, 32'sd453, 32'sd899, 32'sd750,
32'sd1086, 32'sd1793, 32'sd1237, 32'sd733, 32'sd890, 32'sd1371,
32'sd1751, 32'sd1543, 32'sd314, 32'sd847, 32'sd1895, 32'sd1529,
32'sd1773, 32'sd1840, 32'sd580, 32'sd1421, 32'sd245, 32'sd1078,
32'sd367, 32'sd132, 32'sd1390, 32'sd648, 32'sd1053, 32'sd375,
32'sd546, 32'sd1319, 32'sd1288, 32'sd1803, 32'sd439, 32'sd720,
32'sd1095, 32'sd1059, 32'sd1897, 32'sd1033, 32'sd1556, 32'sd1382,
32'sd1106, 32'sd1411, 32'sd164, 32'sd771, 32'sd1366, 32'sd1939,
32'sd378, 32'sd248, 32'sd1987, 32'sd276, 32'sd1173, 32'sd1349,
32'sd1755, 32'sd1640, 32'sd1473, 32'sd1322, 32'sd1503, 32'sd980,
32'sd1675, 32'sd747, 32'sd1151, 32'sd253, 32'sd1499, 32'sd547,
32'sd1883, 32'sd1443, 32'sd1275, 32'sd530, 32'sd714, 32'sd471,
32'sd1266, 32'sd1289, 32'sd582, 32'sd1254, 32'sd1025, 32'sd1814,
32'sd136, 32'sd142, 32'sd1132, 32'sd631, 32'sd1974, 32'sd1217,
32'sd1862, 32'sd1837, 32'sd1360, 32'sd1812, 32'sd446, 32'sd935,
32'sd451, 32'sd450, 32'sd577, 32'sd1250, 32'sd547, 32'sd309,
32'sd1394, 32'sd544, 32'sd1146, 32'sd1944, 32'sd837, 32'sd1498,
32'sd1824, 32'sd1375, 32'sd1493, 32'sd859, 32'sd1737, 32'sd1416,
32'sd1182, 32'sd622, 32'sd1736, 32'sd463, 32'sd245, 32'sd782,
32'sd549, 32'sd786, 32'sd1376, 32'sd871, 32'sd485, 32'sd101,
32'sd1903, 32'sd2000, 32'sd228, 32'sd495, 32'sd580, 32'sd1735,
32'sd483, 32'sd1415, 32'sd182, 32'sd582, 32'sd603, 32'sd905,
32'sd696, 32'sd683, 32'sd389, 32'sd984, 32'sd809, 32'sd430,
32'sd1995, 32'sd461, 32'sd488, 32'sd1694, 32'sd1929, 32'sd662,
32'sd1503, 32'sd1623, 32'sd262, 32'sd1097, 32'sd104, 32'sd537,
32'sd268, 32'sd967, 32'sd864, 32'sd1917, 32'sd583, 32'sd1759,
32'sd1316, 32'sd1864, 32'sd806, 32'sd1018, 32'sd839, 32'sd1210,
32'sd1800, 32'sd598, 32'sd674, 32'sd120, 32'sd1111, 32'sd1424,
32'sd969, 32'sd1967, 32'sd1469, 32'sd1111, 32'sd365, 32'sd1714,
32'sd1871, 32'sd350, 32'sd1829, 32'sd1239, 32'sd1697, 32'sd156,
32'sd391, 32'sd1810, 32'sd1080, 32'sd1689, 32'sd1095, 32'sd849,
32'sd1055, 32'sd405, 32'sd1259, 32'sd348, 32'sd1334, 32'sd1870,
32'sd1284, 32'sd214, 32'sd1009, 32'sd349, 32'sd432, 32'sd1575,
32'sd1267, 32'sd1022, 32'sd943, 32'sd1234, 32'sd1397, 32'sd1721,
32'sd525, 32'sd1208, 32'sd983, 32'sd392, 32'sd1758, 32'sd1725,
32'sd921, 32'sd1910, 32'sd1701, 32'sd1873, 32'sd1901, 32'sd1715,
32'sd1413, 32'sd1037, 32'sd252, 32'sd1660, 32'sd1216, 32'sd859,
32'sd839, 32'sd597, 32'sd823, 32'sd1267, 32'sd311, 32'sd915,
32'sd449, 32'sd782, 32'sd1444, 32'sd1971, 32'sd861, 32'sd998,
32'sd1596, 32'sd254, 32'sd677, 32'sd1842, 32'sd1065, 32'sd1478,
32'sd578, 32'sd1095, 32'sd1897, 32'sd1569, 32'sd613, 32'sd1951,
32'sd844, 32'sd808, 32'sd823, 32'sd769, 32'sd871, 32'sd900,
32'sd862, 32'sd516, 32'sd1305, 32'sd1147, 32'sd1610, 32'sd654,
32'sd1932, 32'sd1024, 32'sd111, 32'sd934, 32'sd272, 32'sd568,
32'sd1850, 32'sd1365, 32'sd469, 32'sd1496, 32'sd1795, 32'sd1022,
32'sd1734, 32'sd1496, 32'sd363, 32'sd356, 32'sd1386, 32'sd1474,
32'sd1656, 32'sd318, 32'sd1177, 32'sd1127, 32'sd1243, 32'sd562,
32'sd153, 32'sd1047, 32'sd1094, 32'sd1409, 32'sd1280, 32'sd1317,
32'sd715, 32'sd1952, 32'sd1960, 32'sd1391, 32'sd1701, 32'sd399,
32'sd559, 32'sd837, 32'sd540, 32'sd196, 32'sd891, 32'sd1179,
32'sd1644, 32'sd578, 32'sd1755, 32'sd675, 32'sd533, 32'sd1965,
32'sd1302, 32'sd361, 32'sd1415, 32'sd824, 32'sd1750, 32'sd1226,
32'sd1929, 32'sd1639, 32'sd1355, 32'sd817, 32'sd1357, 32'sd872,
32'sd903, 32'sd446, 32'sd1434, 32'sd883, 32'sd105, 32'sd1907,
32'sd315, 32'sd1382, 32'sd483, 32'sd1692, 32'sd688, 32'sd202,
32'sd1351, 32'sd548, 32'sd566, 32'sd211, 32'sd146, 32'sd1858,
32'sd524, 32'sd280, 32'sd1647, 32'sd459, 32'sd546, 32'sd1850,
32'sd450, 32'sd159, 32'sd1870, 32'sd1103, 32'sd1494, 32'sd275,
32'sd837, 32'sd1795, 32'sd394, 32'sd1709, 32'sd647, 32'sd1721,
32'sd440, 32'sd273, 32'sd1628, 32'sd896, 32'sd1978, 32'sd1775,
32'sd263, 32'sd988, 32'sd1948, 32'sd490, 32'sd1335, 32'sd1926,
32'sd659, 32'sd677, 32'sd362, 32'sd1727, 32'sd1595, 32'sd1169,
32'sd1695, 32'sd296, 32'sd1430, 32'sd1332, 32'sd839, 32'sd1104,
32'sd458, 32'sd966, 32'sd1715, 32'sd684, 32'sd1273, 32'sd1039,
32'sd1579, 32'sd158, 32'sd1561, 32'sd1663, 32'sd1874, 32'sd866,
32'sd1294, 32'sd629, 32'sd503, 32'sd1874, 32'sd1578, 32'sd1919,
32'sd977, 32'sd701, 32'sd646, 32'sd193, 32'sd1603, 32'sd1633,
32'sd363, 32'sd1278, 32'sd653, 32'sd598, 32'sd1014, 32'sd1552,
32'sd569, 32'sd225, 32'sd1035, 32'sd1028, 32'sd318, 32'sd1920,
32'sd553, 32'sd1416, 32'sd1899, 32'sd347, 32'sd722, 32'sd1925,
32'sd486, 32'sd533, 32'sd1830, 32'sd219, 32'sd827, 32'sd621,
32'sd388, 32'sd1543, 32'sd1421, 32'sd749, 32'sd1090, 32'sd1307,
32'sd407, 32'sd567, 32'sd1249, 32'sd1420, 32'sd1006, 32'sd1513,
32'sd1046, 32'sd1679, 32'sd1481, 32'sd569, 32'sd1851, 32'sd357,
32'sd281, 32'sd1346, 32'sd786, 32'sd687, 32'sd968, 32'sd524,
32'sd398, 32'sd1199, 32'sd578, 32'sd1061, 32'sd1422, 32'sd1388,
32'sd728, 32'sd1825, 32'sd1316, 32'sd637, 32'sd1704, 32'sd626,
32'sd475, 32'sd720, 32'sd1241, 32'sd926, 32'sd1323, 32'sd530,
32'sd534, 32'sd1584, 32'sd600, 32'sd834, 32'sd1065, 32'sd1474,
32'sd847, 32'sd1564, 32'sd1316, 32'sd1445, 32'sd1619, 32'sd522,
32'sd793, 32'sd863, 32'sd633, 32'sd961, 32'sd1357, 32'sd1849,
32'sd443, 32'sd755, 32'sd1863, 32'sd932, 32'sd656, 32'sd1557,
32'sd1147, 32'sd846, 32'sd339, 32'sd1169, 32'sd390, 32'sd1768,
32'sd215, 32'sd242, 32'sd1927, 32'sd231, 32'sd1570, 32'sd1087,
32'sd1871, 32'sd284, 32'sd1406, 32'sd1962, 32'sd1271, 32'sd905,
32'sd1603, 32'sd1489, 32'sd1611, 32'sd165, 32'sd1798, 32'sd1892,
32'sd1401, 32'sd870, 32'sd821, 32'sd555, 32'sd1675, 32'sd972,
32'sd652, 32'sd1136, 32'sd1341, 32'sd1871, 32'sd195, 32'sd224,
32'sd914, 32'sd532, 32'sd378, 32'sd1639, 32'sd1875, 32'sd412,
32'sd217, 32'sd1684, 32'sd141, 32'sd493, 32'sd748, 32'sd231,
32'sd734, 32'sd416, 32'sd197, 32'sd1771, 32'sd1878, 32'sd843,
32'sd1108, 32'sd1188, 32'sd441, 32'sd982, 32'sd1425, 32'sd924,
32'sd1295, 32'sd1279, 32'sd693, 32'sd161, 32'sd1246, 32'sd1424,
32'sd1054, 32'sd286, 32'sd944, 32'sd1982, 32'sd723, 32'sd1462,
32'sd1672, 32'sd1798, 32'sd335, 32'sd1859, 32'sd487, 32'sd634,
32'sd1152, 32'sd992, 32'sd1451, 32'sd1783, 32'sd425, 32'sd260,
32'sd601, 32'sd1806, 32'sd1321, 32'sd1851, 32'sd616, 32'sd1365,
32'sd1863, 32'sd1426, 32'sd1396, 32'sd1632, 32'sd1025, 32'sd476,
32'sd821, 32'sd1907, 32'sd859, 32'sd1203, 32'sd231, 32'sd1193,
32'sd520, 32'sd212, 32'sd1117, 32'sd558, 32'sd1061, 32'sd1764,
32'sd1264, 32'sd1687, 32'sd880, 32'sd1147, 32'sd1092, 32'sd1439,
32'sd1203, 32'sd1135, 32'sd895, 32'sd1889, 32'sd852, 32'sd1701,
32'sd712, 32'sd1942, 32'sd1371, 32'sd460, 32'sd1638, 32'sd1800,
32'sd1622, 32'sd191, 32'sd1424, 32'sd977, 32'sd974, 32'sd560,
32'sd1625, 32'sd1698, 32'sd1774, 32'sd1060, 32'sd1962, 32'sd1365,
32'sd597, 32'sd995, 32'sd1146, 32'sd1354, 32'sd1455, 32'sd119,
32'sd1356, 32'sd1849, 32'sd1208, 32'sd1197, 32'sd521, 32'sd1696,
32'sd1099, 32'sd1516, 32'sd1255, 32'sd597, 32'sd1487, 32'sd126,
32'sd572, 32'sd1077, 32'sd1906, 32'sd930, 32'sd932, 32'sd540,
32'sd1580, 32'sd1015, 32'sd167, 32'sd1401, 32'sd411, 32'sd1265,
32'sd1028, 32'sd889, 32'sd1903, 32'sd1013, 32'sd1075, 32'sd1851,
32'sd1952, 32'sd1000, 32'sd495, 32'sd570, 32'sd1208, 32'sd520,
32'sd1915, 32'sd1906, 32'sd471, 32'sd555, 32'sd328, 32'sd695,
32'sd1579, 32'sd1563, 32'sd1622, 32'sd1918, 32'sd1942, 32'sd1623,
32'sd1698, 32'sd871, 32'sd762, 32'sd1545, 32'sd1739, 32'sd1789,
32'sd792, 32'sd141, 32'sd1027, 32'sd235, 32'sd775, 32'sd1998,
32'sd1133, 32'sd553, 32'sd1734, 32'sd1510, 32'sd992, 32'sd1921,
32'sd1455, 32'sd1777, 32'sd1197, 32'sd595, 32'sd1852, 32'sd112,
32'sd1086, 32'sd1155, 32'sd641, 32'sd165, 32'sd124, 32'sd1680,
32'sd1873, 32'sd704, 32'sd997, 32'sd354, 32'sd437, 32'sd1841,
32'sd1796, 32'sd1143, 32'sd213, 32'sd1253, 32'sd1505, 32'sd1937,
32'sd442, 32'sd1056, 32'sd928, 32'sd970, 32'sd274, 32'sd1863,
32'sd1721, 32'sd1687, 32'sd134, 32'sd129, 32'sd1067, 32'sd106,
32'sd178, 32'sd1169, 32'sd939, 32'sd1768, 32'sd1019, 32'sd1613,
32'sd320, 32'sd776, 32'sd1565, 32'sd1057, 32'sd825, 32'sd1773,
32'sd504, 32'sd340, 32'sd957, 32'sd469, 32'sd1468, 32'sd1010,
32'sd1438, 32'sd1700, 32'sd510, 32'sd974, 32'sd1567, 32'sd1609,
32'sd250, 32'sd1914, 32'sd1526, 32'sd658, 32'sd1675, 32'sd903,
32'sd903, 32'sd1334, 32'sd1496, 32'sd716, 32'sd695, 32'sd1617,
32'sd1517, 32'sd1006, 32'sd1846, 32'sd449, 32'sd172, 32'sd962,
32'sd185, 32'sd935, 32'sd241, 32'sd1471, 32'sd1293, 32'sd1313,
32'sd1925, 32'sd937, 32'sd1995, 32'sd1088, 32'sd1323, 32'sd692,
32'sd1333, 32'sd757, 32'sd814, 32'sd1586, 32'sd1899, 32'sd303,
32'sd1801, 32'sd1697, 32'sd1825, 32'sd1036, 32'sd1683, 32'sd884,
32'sd1021, 32'sd1811, 32'sd793, 32'sd1839, 32'sd218, 32'sd369,
32'sd1612, 32'sd381, 32'sd1798, 32'sd695, 32'sd830, 32'sd1765,
32'sd1235, 32'sd1453, 32'sd1051, 32'sd1221, 32'sd1553, 32'sd887,
32'sd1407, 32'sd994, 32'sd322, 32'sd1371, 32'sd1019, 32'sd672,
32'sd995, 32'sd987, 32'sd425, 32'sd969, 32'sd500, 32'sd246,
32'sd1216, 32'sd1961, 32'sd1989, 32'sd1780, 32'sd1583, 32'sd606,
32'sd424, 32'sd327, 32'sd1048, 32'sd1809, 32'sd794, 32'sd755,
32'sd954, 32'sd853, 32'sd320, 32'sd1355, 32'sd1787, 32'sd1708,
32'sd1853, 32'sd689, 32'sd894, 32'sd354, 32'sd1688, 32'sd162,
32'sd785, 32'sd975, 32'sd158, 32'sd1972, 32'sd216, 32'sd950,
32'sd1257, 32'sd864, 32'sd804, 32'sd602, 32'sd779, 32'sd1492,
32'sd271, 32'sd1239, 32'sd394, 32'sd467, 32'sd1817, 32'sd428,
32'sd1656, 32'sd1522, 32'sd493, 32'sd163, 32'sd842, 32'sd281,
32'sd1290, 32'sd1968, 32'sd785, 32'sd508, 32'sd264, 32'sd680,
32'sd426, 32'sd1146, 32'sd1175, 32'sd734, 32'sd514, 32'sd1283,
32'sd1762, 32'sd1163, 32'sd693, 32'sd1786, 32'sd1611, 32'sd1537,
32'sd974, 32'sd634, 32'sd722, 32'sd1989, 32'sd1280, 32'sd1663,
32'sd1196, 32'sd348, 32'sd1866, 32'sd1386, 32'sd1404, 32'sd880,
32'sd1115, 32'sd254, 32'sd1262, 32'sd856, 32'sd1032, 32'sd567,
32'sd282, 32'sd809, 32'sd1029, 32'sd1191, 32'sd261, 32'sd908,
32'sd674, 32'sd1191, 32'sd1149, 32'sd1505, 32'sd1974, 32'sd1693,
32'sd1831, 32'sd1083, 32'sd1529, 32'sd1831, 32'sd1127, 32'sd819,
32'sd380, 32'sd763, 32'sd1802, 32'sd1822, 32'sd1842, 32'sd706,
32'sd1247, 32'sd350, 32'sd315, 32'sd343, 32'sd928, 32'sd942,
32'sd1541, 32'sd812, 32'sd789, 32'sd1151, 32'sd856, 32'sd974,
32'sd214, 32'sd956, 32'sd1758, 32'sd1565, 32'sd1166, 32'sd232,
32'sd1427, 32'sd1244, 32'sd977, 32'sd1806, 32'sd992, 32'sd1143,
32'sd821, 32'sd165, 32'sd736, 32'sd359, 32'sd1627, 32'sd1303,
32'sd107, 32'sd622, 32'sd454, 32'sd1369, 32'sd139, 32'sd1256,
32'sd490, 32'sd1413, 32'sd1075, 32'sd851, 32'sd611, 32'sd498,
32'sd1079, 32'sd1555, 32'sd663, 32'sd663, 32'sd1620, 32'sd384,
32'sd1207, 32'sd1962, 32'sd1096, 32'sd845, 32'sd1398, 32'sd1799,
32'sd1216, 32'sd1763, 32'sd301, 32'sd956, 32'sd1615, 32'sd960,
32'sd1714, 32'sd1609, 32'sd338, 32'sd1185, 32'sd1875, 32'sd1063,
32'sd782, 32'sd797, 32'sd1584, 32'sd1572, 32'sd627, 32'sd955,
32'sd1417, 32'sd1032, 32'sd1406, 32'sd1433, 32'sd1670, 32'sd1105,
32'sd210, 32'sd758, 32'sd1123, 32'sd716, 32'sd821, 32'sd303,
32'sd379, 32'sd406, 32'sd1825, 32'sd1175, 32'sd1379, 32'sd1201,
32'sd1870, 32'sd1925, 32'sd266, 32'sd304, 32'sd1184, 32'sd1513,
32'sd127, 32'sd107, 32'sd1666, 32'sd1317, 32'sd653, 32'sd363,
32'sd1522, 32'sd117, 32'sd1373, 32'sd1018, 32'sd1827, 32'sd1201,
32'sd781, 32'sd521, 32'sd1773, 32'sd1700, 32'sd634, 32'sd1527,
32'sd1087, 32'sd179, 32'sd1237, 32'sd704, 32'sd1073, 32'sd163,
32'sd1186, 32'sd1764, 32'sd1692, 32'sd391, 32'sd1414, 32'sd1416,
32'sd1767, 32'sd594, 32'sd983, 32'sd1346, 32'sd1346, 32'sd1419,
32'sd967, 32'sd608, 32'sd1704, 32'sd1670, 32'sd168, 32'sd874,
32'sd470, 32'sd849, 32'sd707, 32'sd1068, 32'sd1284, 32'sd585,
32'sd1381, 32'sd468, 32'sd1032, 32'sd1402, 32'sd657, 32'sd638,
32'sd1416, 32'sd1566, 32'sd1519, 32'sd1737, 32'sd1920, 32'sd655,
32'sd962, 32'sd1194, 32'sd308, 32'sd1296, 32'sd341, 32'sd552,
32'sd731, 32'sd1888, 32'sd1353, 32'sd531, 32'sd858, 32'sd789,
32'sd205, 32'sd387, 32'sd117, 32'sd1478, 32'sd1975, 32'sd736,
32'sd1657, 32'sd865, 32'sd1464, 32'sd1336, 32'sd231, 32'sd944,
32'sd778, 32'sd1192, 32'sd510, 32'sd1666, 32'sd596, 32'sd765,
32'sd1067, 32'sd836, 32'sd883, 32'sd116, 32'sd763, 32'sd617,
32'sd1517, 32'sd1197, 32'sd1378, 32'sd1034, 32'sd1767, 32'sd1440,
32'sd1938, 32'sd572, 32'sd1691, 32'sd829, 32'sd399, 32'sd773,
32'sd991, 32'sd530, 32'sd1635, 32'sd1232, 32'sd744, 32'sd237,
32'sd374, 32'sd1498, 32'sd1651, 32'sd1472, 32'sd1937, 32'sd1465,
32'sd895, 32'sd997, 32'sd560, 32'sd1921, 32'sd1037, 32'sd1796,
32'sd322, 32'sd650, 32'sd1529, 32'sd1556, 32'sd1161, 32'sd1840,
32'sd1955, 32'sd204, 32'sd1380, 32'sd802, 32'sd1425, 32'sd770,
32'sd1931, 32'sd1264, 32'sd1110, 32'sd528, 32'sd1625, 32'sd595,
32'sd1641, 32'sd246, 32'sd1528, 32'sd1476, 32'sd902, 32'sd1156,
32'sd1805, 32'sd522, 32'sd916, 32'sd896, 32'sd1016, 32'sd1987,
32'sd276, 32'sd507, 32'sd674, 32'sd1102, 32'sd1162, 32'sd1227,
32'sd716, 32'sd167, 32'sd1044, 32'sd1361, 32'sd1081, 32'sd437,
32'sd530, 32'sd342, 32'sd1569, 32'sd1156, 32'sd1822, 32'sd1413,
32'sd1599, 32'sd1523, 32'sd1825, 32'sd471, 32'sd292, 32'sd662,
32'sd1711, 32'sd102, 32'sd1246, 32'sd1272, 32'sd1823, 32'sd1589,
32'sd1846, 32'sd1013, 32'sd1933, 32'sd1789, 32'sd1204, 32'sd206,
32'sd291, 32'sd1235, 32'sd1302, 32'sd1148, 32'sd1001, 32'sd661,
32'sd628, 32'sd1016, 32'sd529, 32'sd1959, 32'sd1480, 32'sd243,
32'sd1698, 32'sd1334, 32'sd843, 32'sd1419, 32'sd971, 32'sd1118,
32'sd342, 32'sd212, 32'sd1607, 32'sd1561, 32'sd1624, 32'sd1843,
32'sd1198, 32'sd1469, 32'sd250, 32'sd1824, 32'sd226, 32'sd186,
32'sd107, 32'sd1435, 32'sd382, 32'sd1207, 32'sd1821, 32'sd345,
32'sd712, 32'sd1892, 32'sd1806, 32'sd840, 32'sd416, 32'sd1516,
32'sd1642, 32'sd1246, 32'sd1812, 32'sd141, 32'sd485, 32'sd593,
32'sd1374, 32'sd459, 32'sd523, 32'sd810, 32'sd768, 32'sd381,
32'sd313, 32'sd191, 32'sd542, 32'sd219, 32'sd1493, 32'sd351,
32'sd361, 32'sd1624, 32'sd1707, 32'sd1168, 32'sd565, 32'sd1532,
32'sd147, 32'sd351, 32'sd1355, 32'sd138, 32'sd1762, 32'sd124,
32'sd765, 32'sd1414, 32'sd1494, 32'sd1236, 32'sd972, 32'sd962,
32'sd542, 32'sd1585, 32'sd223, 32'sd239, 32'sd268, 32'sd149,
32'sd1045, 32'sd1629, 32'sd568, 32'sd1223, 32'sd984, 32'sd1937,
32'sd372, 32'sd1934, 32'sd1588, 32'sd1518, 32'sd361, 32'sd151,
32'sd1703, 32'sd1637, 32'sd467, 32'sd1656, 32'sd1777, 32'sd1167,
32'sd1619, 32'sd1890, 32'sd1269, 32'sd1707, 32'sd1937, 32'sd1887,
32'sd1711, 32'sd182, 32'sd963, 32'sd706, 32'sd192, 32'sd1631,
32'sd1977, 32'sd1907, 32'sd1556, 32'sd166, 32'sd119, 32'sd1888,
32'sd481, 32'sd295, 32'sd1626, 32'sd712, 32'sd924, 32'sd968,
32'sd245, 32'sd953, 32'sd296, 32'sd1909, 32'sd943, 32'sd542,
32'sd1667, 32'sd693, 32'sd1418, 32'sd1934, 32'sd1263, 32'sd405,
32'sd104, 32'sd1819, 32'sd433, 32'sd998, 32'sd1609, 32'sd829,
32'sd534, 32'sd1605, 32'sd1622, 32'sd1669, 32'sd1654, 32'sd423,
32'sd285, 32'sd1836, 32'sd1836, 32'sd708, 32'sd1808, 32'sd283,
32'sd1953, 32'sd307, 32'sd1960, 32'sd258, 32'sd584, 32'sd136,
32'sd1208, 32'sd290, 32'sd235, 32'sd1976, 32'sd1838, 32'sd1487,
32'sd1598, 32'sd1662, 32'sd1697, 32'sd308, 32'sd1234, 32'sd512,
32'sd1503, 32'sd844, 32'sd794, 32'sd1418, 32'sd1624, 32'sd424,
32'sd873, 32'sd821, 32'sd1328, 32'sd1789, 32'sd1799, 32'sd1378,
32'sd483, 32'sd1992, 32'sd1906, 32'sd1130, 32'sd1776, 32'sd692,
32'sd656, 32'sd1235, 32'sd1326, 32'sd685, 32'sd766, 32'sd795,
32'sd1000, 32'sd1777, 32'sd614, 32'sd1742, 32'sd1036, 32'sd1930,
32'sd1965, 32'sd339, 32'sd678, 32'sd1700, 32'sd1648, 32'sd1721,
32'sd1046, 32'sd351, 32'sd1168, 32'sd549, 32'sd449, 32'sd1927,
32'sd343, 32'sd1438, 32'sd1466, 32'sd1753, 32'sd378, 32'sd262,
32'sd1720, 32'sd132, 32'sd1890, 32'sd847, 32'sd1595, 32'sd1977,
32'sd1371, 32'sd1513, 32'sd1505, 32'sd572, 32'sd1914, 32'sd1513,
32'sd636, 32'sd222, 32'sd574, 32'sd1214, 32'sd391, 32'sd1491,
32'sd1645, 32'sd104, 32'sd1820, 32'sd612, 32'sd159, 32'sd1121,
32'sd1369, 32'sd1304, 32'sd419, 32'sd496, 32'sd1705, 32'sd1964,
32'sd1810, 32'sd356, 32'sd1978, 32'sd1172, 32'sd1169, 32'sd1658,
32'sd1941, 32'sd667, 32'sd1957, 32'sd349, 32'sd942, 32'sd798,
32'sd565, 32'sd428, 32'sd1060, 32'sd1278, 32'sd196, 32'sd1867,
32'sd588, 32'sd1587, 32'sd1085, 32'sd864, 32'sd1714, 32'sd154,
32'sd1533, 32'sd1011, 32'sd1532, 32'sd1898, 32'sd559, 32'sd1569,
32'sd795, 32'sd835, 32'sd1884, 32'sd118, 32'sd1221, 32'sd612,
32'sd437, 32'sd1917, 32'sd392, 32'sd108, 32'sd1313, 32'sd1882,
32'sd1180, 32'sd829, 32'sd836, 32'sd1209, 32'sd639, 32'sd1242,
32'sd567, 32'sd1350, 32'sd1286, 32'sd592, 32'sd708, 32'sd1997,
32'sd1204, 32'sd791, 32'sd1397, 32'sd1246, 32'sd1712, 32'sd437,
32'sd225, 32'sd1796, 32'sd176, 32'sd1094, 32'sd1864, 32'sd1603,
32'sd1388, 32'sd1374, 32'sd835, 32'sd1634, 32'sd335, 32'sd947,
32'sd1926, 32'sd289, 32'sd863, 32'sd1270, 32'sd1434, 32'sd1661,
32'sd775, 32'sd1056, 32'sd1358, 32'sd332, 32'sd1721, 32'sd1911,
32'sd1875, 32'sd1105, 32'sd267, 32'sd1971, 32'sd464, 32'sd146,
32'sd703, 32'sd574, 32'sd1357, 32'sd210, 32'sd222, 32'sd198,
32'sd1142, 32'sd284, 32'sd710, 32'sd1570, 32'sd1097, 32'sd445,
32'sd1620, 32'sd329, 32'sd478, 32'sd164, 32'sd1030, 32'sd1409,
32'sd452, 32'sd1415, 32'sd167, 32'sd801, 32'sd1093, 32'sd713,
32'sd413, 32'sd715, 32'sd1823, 32'sd1600, 32'sd463, 32'sd1354,
32'sd1957, 32'sd350, 32'sd1126, 32'sd212, 32'sd1916, 32'sd569,
32'sd545, 32'sd1035, 32'sd1840, 32'sd664, 32'sd949, 32'sd231,
32'sd1640, 32'sd1714, 32'sd1133, 32'sd1212, 32'sd1660, 32'sd398,
32'sd997, 32'sd862, 32'sd1075, 32'sd163, 32'sd1563, 32'sd1904,
32'sd670, 32'sd361, 32'sd1630, 32'sd362, 32'sd195, 32'sd1195,
32'sd1704, 32'sd1216, 32'sd1153, 32'sd1394, 32'sd701, 32'sd1857,
32'sd529, 32'sd1552, 32'sd1122, 32'sd920, 32'sd814, 32'sd200,
32'sd1007, 32'sd1669, 32'sd1934, 32'sd223, 32'sd548, 32'sd265,
32'sd390, 32'sd1991, 32'sd1228, 32'sd321, 32'sd1380, 32'sd428,
32'sd1431, 32'sd1772, 32'sd225, 32'sd1293, 32'sd1469, 32'sd996,
32'sd162, 32'sd113, 32'sd1088, 32'sd1977, 32'sd951, 32'sd678,
32'sd1440, 32'sd288, 32'sd1980, 32'sd129, 32'sd224, 32'sd1879,
32'sd177, 32'sd980, 32'sd503, 32'sd1043, 32'sd1365, 32'sd825,
32'sd902, 32'sd585, 32'sd1639, 32'sd1676, 32'sd884, 32'sd1790,
32'sd1704, 32'sd692, 32'sd1805, 32'sd812, 32'sd533, 32'sd385,
32'sd1747, 32'sd1740, 32'sd1539, 32'sd1933, 32'sd520, 32'sd1995,
32'sd911, 32'sd1944, 32'sd1731, 32'sd489, 32'sd438, 32'sd1159,
32'sd1522, 32'sd548, 32'sd730, 32'sd410, 32'sd470, 32'sd682,
32'sd1409, 32'sd1291, 32'sd1035, 32'sd1237, 32'sd106, 32'sd893,
32'sd1293, 32'sd643, 32'sd1537, 32'sd399, 32'sd1606, 32'sd135,
32'sd1006, 32'sd965, 32'sd1767, 32'sd1378, 32'sd983, 32'sd341,
32'sd206, 32'sd150, 32'sd290, 32'sd948, 32'sd121, 32'sd1250,
32'sd888, 32'sd980, 32'sd1324, 32'sd424, 32'sd1112, 32'sd1706,
32'sd777, 32'sd208, 32'sd338, 32'sd421, 32'sd179, 32'sd1016,
32'sd968, 32'sd1546, 32'sd477, 32'sd984, 32'sd1678, 32'sd597,
32'sd173, 32'sd556, 32'sd170, 32'sd745, 32'sd1018, 32'sd1421,
32'sd1485, 32'sd316, 32'sd1720, 32'sd1590, 32'sd1055, 32'sd579,
32'sd916, 32'sd1275, 32'sd1275, 32'sd1494, 32'sd584, 32'sd559,
32'sd1547, 32'sd344, 32'sd1790, 32'sd1981, 32'sd1416, 32'sd1399,
32'sd1897, 32'sd1785, 32'sd1862, 32'sd1314, 32'sd471, 32'sd598,
32'sd287, 32'sd579, 32'sd1475, 32'sd1657, 32'sd1926, 32'sd1992,
32'sd1151, 32'sd1933, 32'sd1930, 32'sd1881, 32'sd1821, 32'sd152,
32'sd1587, 32'sd101, 32'sd1649, 32'sd418, 32'sd1110, 32'sd707,
32'sd652, 32'sd1557, 32'sd1398, 32'sd514, 32'sd1798, 32'sd1753,
32'sd1490, 32'sd692, 32'sd1986, 32'sd1848, 32'sd1061, 32'sd516,
32'sd262, 32'sd428, 32'sd331, 32'sd1662, 32'sd1017, 32'sd614,
32'sd955, 32'sd772, 32'sd104, 32'sd1361, 32'sd1170, 32'sd638,
32'sd1089, 32'sd651, 32'sd1359, 32'sd1546, 32'sd568, 32'sd1128,
32'sd399, 32'sd472, 32'sd1664, 32'sd1643, 32'sd735, 32'sd1049,
32'sd1179, 32'sd198, 32'sd1686, 32'sd1746, 32'sd422, 32'sd1483,
32'sd293, 32'sd1709, 32'sd1929, 32'sd1265, 32'sd916, 32'sd237,
32'sd1911, 32'sd1574, 32'sd1657, 32'sd1286, 32'sd166, 32'sd1329,
32'sd141, 32'sd1552, 32'sd1379, 32'sd1386, 32'sd659, 32'sd720,
32'sd1335, 32'sd318, 32'sd406, 32'sd865, 32'sd425, 32'sd1144,
32'sd768, 32'sd876, 32'sd727, 32'sd1710, 32'sd796, 32'sd1043,
32'sd495, 32'sd1404, 32'sd894, 32'sd1175, 32'sd1831, 32'sd1076,
32'sd1983, 32'sd1434, 32'sd1204, 32'sd280, 32'sd543, 32'sd1366,
32'sd1641, 32'sd369, 32'sd1097, 32'sd1275, 32'sd254, 32'sd1552,
32'sd738, 32'sd1108, 32'sd1807, 32'sd1943, 32'sd1278, 32'sd624,
32'sd1473, 32'sd1240, 32'sd1187, 32'sd1180, 32'sd1459, 32'sd1607,
32'sd1978, 32'sd316, 32'sd1422, 32'sd998, 32'sd1140, 32'sd1669,
32'sd1281, 32'sd1500, 32'sd777, 32'sd1468, 32'sd1110, 32'sd1565,
32'sd170, 32'sd432, 32'sd1040, 32'sd997, 32'sd115, 32'sd1108,
32'sd1966, 32'sd1112, 32'sd464, 32'sd270, 32'sd1990, 32'sd898,
32'sd1129, 32'sd1016, 32'sd1076, 32'sd863, 32'sd1235, 32'sd1819,
32'sd1306, 32'sd1222, 32'sd462, 32'sd1270, 32'sd942, 32'sd1599,
32'sd868, 32'sd401, 32'sd125, 32'sd1328, 32'sd420, 32'sd479,
32'sd1570, 32'sd1401, 32'sd928, 32'sd998, 32'sd397, 32'sd265,
32'sd977, 32'sd1573, 32'sd926, 32'sd1900, 32'sd134, 32'sd996,
32'sd1556, 32'sd664, 32'sd804, 32'sd805, 32'sd256, 32'sd1268,
32'sd806, 32'sd199, 32'sd1125, 32'sd1432, 32'sd1625, 32'sd379,
32'sd1375, 32'sd639, 32'sd621, 32'sd1509, 32'sd580, 32'sd1465,
32'sd316, 32'sd358, 32'sd112, 32'sd314, 32'sd1416, 32'sd1332,
32'sd1003, 32'sd1678, 32'sd778, 32'sd840, 32'sd1970, 32'sd711,
32'sd1613, 32'sd1046, 32'sd1320, 32'sd297, 32'sd1702, 32'sd1869,
32'sd907, 32'sd1568, 32'sd1424, 32'sd1817, 32'sd1646, 32'sd1810,
32'sd1687, 32'sd1180, 32'sd876, 32'sd1177, 32'sd1244, 32'sd1631,
32'sd332, 32'sd1604, 32'sd1350, 32'sd1262, 32'sd1602, 32'sd1015,
32'sd1429, 32'sd738, 32'sd592, 32'sd1648, 32'sd1351, 32'sd1846,
32'sd1584, 32'sd845, 32'sd364, 32'sd245, 32'sd437, 32'sd460,
32'sd165, 32'sd770, 32'sd396, 32'sd598, 32'sd1124, 32'sd1980,
32'sd1449, 32'sd357, 32'sd1000, 32'sd591, 32'sd645, 32'sd1115,
32'sd1892, 32'sd504, 32'sd958, 32'sd106, 32'sd281, 32'sd1196,
32'sd314, 32'sd313, 32'sd342, 32'sd1523, 32'sd633, 32'sd266,
32'sd875, 32'sd1465, 32'sd1060, 32'sd578, 32'sd1949, 32'sd151,
32'sd226, 32'sd1083, 32'sd1790, 32'sd1074, 32'sd317, 32'sd192,
32'sd1499, 32'sd327, 32'sd1529, 32'sd134, 32'sd707, 32'sd1264,
32'sd1543, 32'sd638, 32'sd1760, 32'sd850, 32'sd1539, 32'sd460,
32'sd1477, 32'sd601, 32'sd1103, 32'sd1083, 32'sd1969, 32'sd1557,
32'sd780, 32'sd1580, 32'sd1911, 32'sd1194, 32'sd1237, 32'sd946,
32'sd1779, 32'sd1100, 32'sd1421, 32'sd831, 32'sd1200, 32'sd1604,
32'sd287, 32'sd1660, 32'sd1001, 32'sd886, 32'sd654, 32'sd1694,
32'sd1429, 32'sd347, 32'sd1835, 32'sd523, 32'sd1098, 32'sd455,
32'sd335, 32'sd1166, 32'sd1320, 32'sd1130, 32'sd865, 32'sd676,
32'sd190, 32'sd628, 32'sd420, 32'sd1392, 32'sd1052, 32'sd920,
32'sd1230, 32'sd717, 32'sd1453, 32'sd1129, 32'sd109, 32'sd941,
32'sd1057, 32'sd1996, 32'sd1904, 32'sd1927, 32'sd886, 32'sd1323,
32'sd696, 32'sd1515, 32'sd1707, 32'sd811, 32'sd1878, 32'sd1448,
32'sd1978, 32'sd1325, 32'sd1997, 32'sd1100, 32'sd1228, 32'sd1045,
32'sd1478, 32'sd713, 32'sd713, 32'sd594, 32'sd1830, 32'sd920,
32'sd1758, 32'sd1830, 32'sd1284, 32'sd1083, 32'sd627, 32'sd1946,
32'sd980, 32'sd387, 32'sd1646, 32'sd911, 32'sd1591, 32'sd256,
32'sd1008, 32'sd101, 32'sd749, 32'sd612, 32'sd519, 32'sd1689,
32'sd1725, 32'sd779, 32'sd455, 32'sd1896, 32'sd1894, 32'sd1799,
32'sd917, 32'sd363, 32'sd1163, 32'sd1566, 32'sd111, 32'sd1545,
32'sd1145, 32'sd439, 32'sd783, 32'sd991, 32'sd683, 32'sd221,
32'sd1714, 32'sd1506, 32'sd1829, 32'sd1295, 32'sd861, 32'sd1825,
32'sd712, 32'sd859, 32'sd1404, 32'sd1340, 32'sd1289, 32'sd630,
32'sd1164, 32'sd934, 32'sd311, 32'sd1942, 32'sd1283, 32'sd541,
32'sd1334, 32'sd1580, 32'sd1966, 32'sd406, 32'sd1929, 32'sd583,
32'sd476, 32'sd1711, 32'sd793, 32'sd985, 32'sd162, 32'sd592,
32'sd815, 32'sd1572, 32'sd1215, 32'sd389, 32'sd1205, 32'sd1734,
32'sd1354, 32'sd1364, 32'sd873, 32'sd835, 32'sd1808, 32'sd1892,
32'sd861, 32'sd565, 32'sd732, 32'sd613, 32'sd363, 32'sd1492,
32'sd1975, 32'sd684, 32'sd886, 32'sd1471, 32'sd1032, 32'sd810,
32'sd529, 32'sd182, 32'sd841, 32'sd1157, 32'sd1004, 32'sd300,
32'sd1527, 32'sd1730, 32'sd1218, 32'sd1796, 32'sd1469, 32'sd1131,
32'sd1857, 32'sd624, 32'sd1481, 32'sd978, 32'sd1514, 32'sd1863,
32'sd805, 32'sd1277, 32'sd496, 32'sd1976, 32'sd1100, 32'sd919,
32'sd330, 32'sd794, 32'sd522, 32'sd897, 32'sd1985, 32'sd471,
32'sd1018, 32'sd1412, 32'sd1533, 32'sd1087, 32'sd1877, 32'sd1561,
32'sd101, 32'sd867, 32'sd1807, 32'sd382, 32'sd1810, 32'sd1435,
32'sd1844, 32'sd1581, 32'sd103, 32'sd688, 32'sd151, 32'sd226,
32'sd1618, 32'sd161, 32'sd1300, 32'sd127, 32'sd1233, 32'sd1362,
32'sd457, 32'sd1791, 32'sd760, 32'sd232, 32'sd786, 32'sd1448,
32'sd854, 32'sd869, 32'sd415, 32'sd858, 32'sd352, 32'sd1573,
32'sd1880, 32'sd826, 32'sd1019, 32'sd142, 32'sd638, 32'sd1469,
32'sd723, 32'sd1389, 32'sd1359, 32'sd1436, 32'sd1217, 32'sd966,
32'sd145, 32'sd1983, 32'sd1302, 32'sd1394, 32'sd602, 32'sd991,
32'sd1560, 32'sd1585, 32'sd572, 32'sd165, 32'sd189, 32'sd606,
32'sd1483, 32'sd1121, 32'sd1182, 32'sd1905, 32'sd1264, 32'sd1837,
32'sd1104, 32'sd1786, 32'sd160, 32'sd1229, 32'sd1003, 32'sd1605,
32'sd724, 32'sd1482, 32'sd1446, 32'sd1451, 32'sd1706, 32'sd1177,
32'sd1116, 32'sd118, 32'sd760, 32'sd139, 32'sd1533, 32'sd1145,
32'sd1347, 32'sd661, 32'sd1227, 32'sd1432, 32'sd1322, 32'sd1662,
32'sd288, 32'sd1448, 32'sd299, 32'sd1863, 32'sd807, 32'sd1812,
32'sd1328, 32'sd230, 32'sd792, 32'sd941, 32'sd560, 32'sd1662,
32'sd1342, 32'sd764, 32'sd572, 32'sd1397, 32'sd702, 32'sd1711,
32'sd1262, 32'sd1616, 32'sd314, 32'sd719, 32'sd1566, 32'sd152,
32'sd1765, 32'sd376, 32'sd739, 32'sd559, 32'sd1764, 32'sd1157,
32'sd726, 32'sd225, 32'sd1841, 32'sd737, 32'sd416, 32'sd738,
32'sd1956, 32'sd1451, 32'sd1595, 32'sd786, 32'sd269, 32'sd579,
32'sd427, 32'sd1129, 32'sd1886, 32'sd1757, 32'sd1146, 32'sd485,
32'sd988, 32'sd1578, 32'sd841, 32'sd125, 32'sd792, 32'sd1526,
32'sd1657, 32'sd1460, 32'sd1010, 32'sd1874, 32'sd1809, 32'sd898,
32'sd1517, 32'sd833, 32'sd1321, 32'sd1875, 32'sd900, 32'sd458,
32'sd1900, 32'sd1453, 32'sd1880, 32'sd262, 32'sd242, 32'sd276,
32'sd442, 32'sd2000, 32'sd1354, 32'sd1664, 32'sd888, 32'sd266,
32'sd271, 32'sd1454, 32'sd1640, 32'sd123, 32'sd1291, 32'sd867,
32'sd1351, 32'sd642, 32'sd1596, 32'sd1563, 32'sd322, 32'sd1888,
32'sd1137, 32'sd933, 32'sd1249, 32'sd1383, 32'sd1598, 32'sd665,
32'sd563, 32'sd1139, 32'sd1527, 32'sd1185, 32'sd1317, 32'sd207,
32'sd1315, 32'sd1831, 32'sd1242, 32'sd1659, 32'sd932, 32'sd216,
32'sd1069, 32'sd942, 32'sd957, 32'sd1879, 32'sd1477, 32'sd1564,
32'sd1741, 32'sd245, 32'sd1469, 32'sd832, 32'sd1248, 32'sd1734,
32'sd298, 32'sd940, 32'sd1976, 32'sd821, 32'sd424, 32'sd642,
32'sd1402, 32'sd273, 32'sd293, 32'sd1292, 32'sd567, 32'sd180,
32'sd1342, 32'sd826, 32'sd1781, 32'sd935, 32'sd1196, 32'sd1308,
32'sd140, 32'sd1553, 32'sd1617, 32'sd960, 32'sd1436, 32'sd1341,
32'sd563, 32'sd1012, 32'sd993, 32'sd1793, 32'sd1388, 32'sd1178,
32'sd449, 32'sd377, 32'sd1809, 32'sd1639, 32'sd469, 32'sd1801,
32'sd225, 32'sd1480, 32'sd957, 32'sd1390, 32'sd800, 32'sd1074,
32'sd1960, 32'sd1247, 32'sd1820, 32'sd304, 32'sd657, 32'sd105,
32'sd1240, 32'sd1386, 32'sd1915, 32'sd472, 32'sd139, 32'sd455,
32'sd1069, 32'sd798, 32'sd942, 32'sd971, 32'sd283, 32'sd1577,
32'sd1167, 32'sd682, 32'sd1341, 32'sd265, 32'sd720, 32'sd1385,
32'sd192, 32'sd886, 32'sd529, 32'sd724, 32'sd438, 32'sd1406,
32'sd887, 32'sd495, 32'sd1818, 32'sd1585, 32'sd1489, 32'sd419,
32'sd812, 32'sd423, 32'sd815, 32'sd1949, 32'sd520, 32'sd182,
32'sd531, 32'sd1769, 32'sd410, 32'sd1350, 32'sd1718, 32'sd1049,
32'sd403, 32'sd1272, 32'sd1572, 32'sd1550, 32'sd1467, 32'sd739,
32'sd1270, 32'sd959, 32'sd148, 32'sd1328, 32'sd221, 32'sd872,
32'sd1612, 32'sd918, 32'sd801, 32'sd687, 32'sd115, 32'sd1092,
32'sd142, 32'sd1174, 32'sd1515, 32'sd522, 32'sd1603, 32'sd856,
32'sd1449, 32'sd1877, 32'sd971, 32'sd157, 32'sd1324, 32'sd459,
32'sd847, 32'sd645, 32'sd1933, 32'sd317, 32'sd554, 32'sd1628,
32'sd448, 32'sd144, 32'sd1604, 32'sd611, 32'sd1925, 32'sd286,
32'sd996, 32'sd1924, 32'sd1820, 32'sd946, 32'sd1075, 32'sd263,
32'sd1402, 32'sd1382, 32'sd300, 32'sd861, 32'sd456, 32'sd1242,
32'sd1815, 32'sd876, 32'sd442, 32'sd226, 32'sd155, 32'sd1303,
32'sd455, 32'sd1847, 32'sd1766, 32'sd254, 32'sd1970, 32'sd413,
32'sd274, 32'sd1749, 32'sd677, 32'sd1760, 32'sd1370, 32'sd565,
32'sd706, 32'sd1343, 32'sd1525, 32'sd1664, 32'sd194, 32'sd1151,
32'sd738, 32'sd1862, 32'sd836, 32'sd1701, 32'sd172, 32'sd1976,
32'sd976, 32'sd1212, 32'sd488, 32'sd1379, 32'sd1840, 32'sd1845,
32'sd704, 32'sd268, 32'sd911, 32'sd1965, 32'sd988, 32'sd161,
32'sd1521, 32'sd445, 32'sd1482, 32'sd351, 32'sd1916, 32'sd1164,
32'sd799, 32'sd191, 32'sd304, 32'sd1423, 32'sd718, 32'sd704,
32'sd1323, 32'sd132, 32'sd984, 32'sd799, 32'sd1779, 32'sd1118,
32'sd922, 32'sd132, 32'sd980, 32'sd393, 32'sd1836, 32'sd1140,
32'sd166, 32'sd1428, 32'sd1115, 32'sd1927, 32'sd1999, 32'sd225,
32'sd1350, 32'sd1957, 32'sd1201, 32'sd953, 32'sd335, 32'sd847,
32'sd295, 32'sd1437, 32'sd288, 32'sd142, 32'sd513, 32'sd1385,
32'sd603, 32'sd1084, 32'sd323, 32'sd1624, 32'sd1831, 32'sd1413,
32'sd1860, 32'sd163, 32'sd140, 32'sd1137, 32'sd1789, 32'sd173,
32'sd352, 32'sd1406, 32'sd892, 32'sd616, 32'sd1013, 32'sd807,
32'sd711, 32'sd1783, 32'sd822, 32'sd1230, 32'sd938, 32'sd1308,
32'sd1176, 32'sd815, 32'sd195, 32'sd383, 32'sd1731, 32'sd740,
32'sd640, 32'sd1005, 32'sd846, 32'sd1013, 32'sd773, 32'sd773,
32'sd1961, 32'sd1470, 32'sd432, 32'sd1010, 32'sd1061, 32'sd1012,
32'sd585, 32'sd1453, 32'sd248, 32'sd325, 32'sd1730, 32'sd723,
32'sd1364, 32'sd1253, 32'sd1408, 32'sd141, 32'sd870, 32'sd225,
32'sd1832, 32'sd1314, 32'sd1358, 32'sd1553, 32'sd940, 32'sd156,
32'sd1517, 32'sd1007, 32'sd1285, 32'sd1438, 32'sd476, 32'sd856,
32'sd1149, 32'sd778, 32'sd130, 32'sd1505, 32'sd1320, 32'sd118,
32'sd1833, 32'sd1133, 32'sd608, 32'sd1267, 32'sd1422, 32'sd1850,
32'sd1493, 32'sd1817, 32'sd949, 32'sd1445, 32'sd1732, 32'sd192,
32'sd196, 32'sd1829, 32'sd128, 32'sd295, 32'sd210, 32'sd1755,
32'sd665, 32'sd411, 32'sd1051, 32'sd698, 32'sd511, 32'sd798,
32'sd1807, 32'sd126, 32'sd1771, 32'sd1146, 32'sd1463, 32'sd330,
32'sd1283, 32'sd1052, 32'sd1879, 32'sd1291, 32'sd600, 32'sd986,
32'sd1601, 32'sd150, 32'sd457, 32'sd1790, 32'sd1068, 32'sd1477,
32'sd1738, 32'sd1382, 32'sd564, 32'sd661, 32'sd1564, 32'sd1822,
32'sd313, 32'sd893, 32'sd1204, 32'sd1190, 32'sd1427, 32'sd882,
32'sd801, 32'sd402, 32'sd1479, 32'sd1093, 32'sd1144, 32'sd186,
32'sd1508, 32'sd1678, 32'sd1247, 32'sd922, 32'sd547, 32'sd296,
32'sd1783, 32'sd1915, 32'sd1893, 32'sd589, 32'sd605, 32'sd365,
32'sd463, 32'sd1417, 32'sd1179, 32'sd1830, 32'sd928, 32'sd613,
32'sd1385, 32'sd1110, 32'sd1926, 32'sd1634, 32'sd1561, 32'sd492,
32'sd814, 32'sd1474, 32'sd1877, 32'sd1009, 32'sd218, 32'sd1626,
32'sd368, 32'sd376, 32'sd1458, 32'sd1000, 32'sd539, 32'sd1180,
32'sd386, 32'sd1118, 32'sd1935, 32'sd753, 32'sd1794, 32'sd685,
32'sd1101, 32'sd891, 32'sd355, 32'sd1954, 32'sd1975, 32'sd1370,
32'sd691, 32'sd1656, 32'sd728, 32'sd1687, 32'sd1535, 32'sd1706,
32'sd291, 32'sd316, 32'sd138, 32'sd1964, 32'sd1705, 32'sd1043,
32'sd1314, 32'sd1754, 32'sd443, 32'sd1036, 32'sd1614, 32'sd1586,
32'sd1515, 32'sd495, 32'sd903, 32'sd426, 32'sd409, 32'sd392,
32'sd1123, 32'sd421, 32'sd1520, 32'sd1103, 32'sd895, 32'sd681,
32'sd400, 32'sd999, 32'sd925, 32'sd1573, 32'sd103, 32'sd432,
32'sd1226, 32'sd259, 32'sd845, 32'sd1634, 32'sd1122, 32'sd141,
32'sd287, 32'sd280, 32'sd109, 32'sd1719, 32'sd201, 32'sd339,
32'sd1736, 32'sd1079, 32'sd537, 32'sd1049, 32'sd974, 32'sd1512,
32'sd946, 32'sd463, 32'sd1214, 32'sd231, 32'sd925, 32'sd623,
32'sd1123, 32'sd392, 32'sd501, 32'sd1485, 32'sd549, 32'sd1855,
32'sd1118, 32'sd867, 32'sd1826, 32'sd1645, 32'sd567, 32'sd1312,
32'sd852, 32'sd1708, 32'sd734, 32'sd1796, 32'sd835, 32'sd883,
32'sd1621, 32'sd1437, 32'sd190, 32'sd663, 32'sd545, 32'sd1502,
32'sd726, 32'sd922, 32'sd1269, 32'sd1025, 32'sd905, 32'sd1563,
32'sd431, 32'sd1730, 32'sd1991, 32'sd478, 32'sd1529, 32'sd705,
32'sd286, 32'sd181, 32'sd305, 32'sd700, 32'sd1846, 32'sd1902,
32'sd1537, 32'sd709, 32'sd601, 32'sd1755, 32'sd1476, 32'sd1322,
32'sd1584, 32'sd1333, 32'sd1521, 32'sd1410, 32'sd555, 32'sd1257,
32'sd631, 32'sd366, 32'sd703, 32'sd706, 32'sd1211, 32'sd1260,
32'sd1232, 32'sd860, 32'sd1411, 32'sd1322, 32'sd1601, 32'sd225,
32'sd993, 32'sd391, 32'sd840, 32'sd402, 32'sd974, 32'sd196,
32'sd165, 32'sd704, 32'sd709, 32'sd271, 32'sd734, 32'sd1662,
32'sd1126, 32'sd669, 32'sd1428, 32'sd1880, 32'sd924, 32'sd583,
32'sd1407, 32'sd594, 32'sd1355, 32'sd1491, 32'sd894, 32'sd1751,
32'sd153, 32'sd1548, 32'sd728, 32'sd320, 32'sd615, 32'sd1714,
32'sd1569, 32'sd1550, 32'sd704, 32'sd438, 32'sd1344, 32'sd444,
32'sd532, 32'sd870, 32'sd1800, 32'sd272, 32'sd604, 32'sd1329,
32'sd842, 32'sd646, 32'sd1200, 32'sd1747, 32'sd851, 32'sd1674,
32'sd685, 32'sd1185, 32'sd225, 32'sd1867, 32'sd1113, 32'sd1778,
32'sd1429, 32'sd1258, 32'sd1649, 32'sd788, 32'sd272, 32'sd1152,
32'sd568, 32'sd246, 32'sd1410, 32'sd1941, 32'sd1803, 32'sd961,
32'sd985, 32'sd539, 32'sd405, 32'sd570, 32'sd721, 32'sd1687,
32'sd1286, 32'sd1925, 32'sd1779, 32'sd1054, 32'sd962, 32'sd1453,
32'sd1423, 32'sd639, 32'sd1298, 32'sd1069, 32'sd1460, 32'sd827,
32'sd1970, 32'sd843, 32'sd610, 32'sd514, 32'sd834, 32'sd1201,
32'sd1181, 32'sd1716, 32'sd1736, 32'sd1694, 32'sd1980, 32'sd1752,
32'sd943, 32'sd1536, 32'sd1794, 32'sd875, 32'sd1418, 32'sd1238,
32'sd719, 32'sd742, 32'sd1391, 32'sd1778, 32'sd446, 32'sd1805,
32'sd1453, 32'sd1048, 32'sd797, 32'sd1337, 32'sd1218, 32'sd499,
32'sd1483, 32'sd1537, 32'sd709, 32'sd1843, 32'sd1815, 32'sd1366,
32'sd212, 32'sd158, 32'sd534, 32'sd1007, 32'sd1005, 32'sd1713,
32'sd1441, 32'sd553, 32'sd1597, 32'sd148, 32'sd1413, 32'sd1930,
32'sd1174, 32'sd1319, 32'sd1676, 32'sd1898, 32'sd110, 32'sd1186,
32'sd1347, 32'sd1675, 32'sd1257, 32'sd1879, 32'sd1978, 32'sd1977,
32'sd1428, 32'sd364, 32'sd1653, 32'sd1701, 32'sd895, 32'sd1239,
32'sd1664, 32'sd1368, 32'sd667, 32'sd1029, 32'sd1312, 32'sd523,
32'sd1341, 32'sd1833, 32'sd1314, 32'sd1157, 32'sd198, 32'sd153,
32'sd1261, 32'sd1695, 32'sd373, 32'sd1070, 32'sd1058, 32'sd1744,
32'sd1051, 32'sd251, 32'sd229, 32'sd250, 32'sd448, 32'sd177,
32'sd1315, 32'sd921, 32'sd1850, 32'sd439, 32'sd1380, 32'sd175,
32'sd1900, 32'sd286, 32'sd841, 32'sd232, 32'sd1111, 32'sd230,
32'sd129, 32'sd1999, 32'sd1563, 32'sd141, 32'sd247, 32'sd1758,
32'sd543, 32'sd387, 32'sd1991, 32'sd1622, 32'sd645, 32'sd1570,
32'sd1837, 32'sd1249, 32'sd1636, 32'sd1028, 32'sd154, 32'sd517,
32'sd1038, 32'sd635, 32'sd265, 32'sd1824, 32'sd413, 32'sd1875,
32'sd1258, 32'sd196, 32'sd384, 32'sd1990, 32'sd1231, 32'sd477,
32'sd293, 32'sd1054, 32'sd211, 32'sd727, 32'sd1095, 32'sd516,
32'sd785, 32'sd231, 32'sd1438, 32'sd1971, 32'sd551, 32'sd1176,
32'sd1385, 32'sd1429, 32'sd293, 32'sd956, 32'sd1592, 32'sd1801,
32'sd949, 32'sd1327, 32'sd1006, 32'sd769, 32'sd425, 32'sd1303,
32'sd609, 32'sd1051, 32'sd1010, 32'sd1074, 32'sd772, 32'sd729,
32'sd474, 32'sd808, 32'sd732, 32'sd1929, 32'sd1236, 32'sd836,
32'sd425, 32'sd787, 32'sd1677, 32'sd187, 32'sd778, 32'sd490,
32'sd706, 32'sd1813, 32'sd519, 32'sd1798, 32'sd153, 32'sd1037,
32'sd1874, 32'sd203, 32'sd1868, 32'sd1649, 32'sd1407, 32'sd642,
32'sd1459, 32'sd1473, 32'sd309, 32'sd208, 32'sd1686, 32'sd1712,
32'sd301, 32'sd686, 32'sd406, 32'sd672, 32'sd1127, 32'sd609,
32'sd1008, 32'sd863, 32'sd107, 32'sd774, 32'sd154, 32'sd1984,
32'sd1981, 32'sd1937, 32'sd657, 32'sd1921, 32'sd1009, 32'sd630,
32'sd915, 32'sd1322, 32'sd1714, 32'sd664, 32'sd1493, 32'sd733,
32'sd746, 32'sd1030, 32'sd1227, 32'sd184, 32'sd1529, 32'sd1617,
32'sd1468, 32'sd1039, 32'sd774, 32'sd581, 32'sd815, 32'sd231,
32'sd1191, 32'sd605, 32'sd1827, 32'sd1611, 32'sd565, 32'sd476,
32'sd456, 32'sd530, 32'sd772, 32'sd1809, 32'sd1703, 32'sd383,
32'sd1384, 32'sd1409, 32'sd276, 32'sd1693, 32'sd1945, 32'sd1279,
32'sd1649, 32'sd1344, 32'sd904, 32'sd889, 32'sd1147, 32'sd632,
32'sd383, 32'sd1911, 32'sd300, 32'sd289, 32'sd1360, 32'sd1437,
32'sd1473, 32'sd479, 32'sd1988, 32'sd1492, 32'sd1964, 32'sd1082,
32'sd1013, 32'sd1574, 32'sd767, 32'sd1506, 32'sd469, 32'sd806,
32'sd685, 32'sd650, 32'sd390, 32'sd217, 32'sd898, 32'sd1252,
32'sd1364, 32'sd1891, 32'sd1222, 32'sd1610, 32'sd1120, 32'sd1991,
32'sd1571, 32'sd1015, 32'sd1645, 32'sd554, 32'sd1057, 32'sd264,
32'sd1458, 32'sd484, 32'sd968, 32'sd1084, 32'sd1976, 32'sd485,
32'sd120, 32'sd1897, 32'sd581, 32'sd987, 32'sd1701, 32'sd1129,
32'sd401, 32'sd1468, 32'sd1275, 32'sd919, 32'sd760, 32'sd953,
32'sd295, 32'sd1032, 32'sd1564, 32'sd766, 32'sd588, 32'sd1335,
32'sd620, 32'sd377, 32'sd1217, 32'sd1938, 32'sd1782, 32'sd552,
32'sd816, 32'sd1588, 32'sd445, 32'sd1210, 32'sd248, 32'sd940,
32'sd245, 32'sd780, 32'sd735, 32'sd567, 32'sd917, 32'sd1467,
32'sd971, 32'sd1101, 32'sd324, 32'sd1057, 32'sd1473, 32'sd164,
32'sd1444, 32'sd703, 32'sd1590, 32'sd751, 32'sd1101, 32'sd130,
32'sd448, 32'sd1545, 32'sd1586, 32'sd795, 32'sd802, 32'sd998,
32'sd450, 32'sd929, 32'sd480, 32'sd1245, 32'sd604, 32'sd270,
32'sd986, 32'sd450, 32'sd207, 32'sd262, 32'sd1710, 32'sd1948,
32'sd1369, 32'sd1262, 32'sd1941, 32'sd689, 32'sd1354, 32'sd1034,
32'sd882, 32'sd711, 32'sd1875, 32'sd756, 32'sd742, 32'sd1771,
32'sd1293, 32'sd587, 32'sd684, 32'sd424, 32'sd603, 32'sd638,
32'sd315, 32'sd1506, 32'sd1251, 32'sd1653, 32'sd881, 32'sd1261,
32'sd1051, 32'sd928, 32'sd1260, 32'sd1803, 32'sd1359, 32'sd928,
32'sd343, 32'sd209, 32'sd1335, 32'sd447, 32'sd1942, 32'sd1847,
32'sd1227, 32'sd1869, 32'sd1690, 32'sd835, 32'sd598, 32'sd1654,
32'sd836, 32'sd590, 32'sd1123, 32'sd1432, 32'sd1889, 32'sd403,
32'sd1825, 32'sd1660, 32'sd1151, 32'sd162, 32'sd1609, 32'sd1190,
32'sd584, 32'sd1372, 32'sd1436, 32'sd1837, 32'sd1559, 32'sd1990,
32'sd395, 32'sd609, 32'sd1363, 32'sd1468, 32'sd1276, 32'sd811,
32'sd103, 32'sd1393, 32'sd184, 32'sd1094, 32'sd529, 32'sd1496,
32'sd1074, 32'sd1285, 32'sd698, 32'sd866, 32'sd1601, 32'sd1770,
32'sd380, 32'sd1115, 32'sd392, 32'sd538, 32'sd864, 32'sd1090,
32'sd1844, 32'sd1956, 32'sd718, 32'sd1710, 32'sd1783, 32'sd207,
32'sd1969, 32'sd932, 32'sd1053, 32'sd1643, 32'sd1948, 32'sd1498,
32'sd205, 32'sd1500, 32'sd1954, 32'sd472, 32'sd1066, 32'sd319,
32'sd1310, 32'sd623, 32'sd587, 32'sd269, 32'sd178, 32'sd1151,
32'sd494, 32'sd1549, 32'sd1262, 32'sd1268, 32'sd1087, 32'sd1872,
32'sd516, 32'sd960, 32'sd1745, 32'sd268, 32'sd1955, 32'sd1545,
32'sd697, 32'sd507, 32'sd1062, 32'sd567, 32'sd830, 32'sd449,
32'sd210, 32'sd773, 32'sd979, 32'sd916, 32'sd322, 32'sd403,
32'sd870, 32'sd718, 32'sd584, 32'sd1671, 32'sd830, 32'sd848,
32'sd251, 32'sd606, 32'sd1428, 32'sd433, 32'sd1407, 32'sd691,
32'sd149, 32'sd618, 32'sd110, 32'sd826, 32'sd413, 32'sd1732,
32'sd1136, 32'sd749, 32'sd505, 32'sd1015, 32'sd1315, 32'sd922,
32'sd614, 32'sd1756, 32'sd1100, 32'sd397, 32'sd1563, 32'sd363,
32'sd1357, 32'sd987, 32'sd1593, 32'sd1759, 32'sd1662, 32'sd1915,
32'sd803, 32'sd1642, 32'sd693, 32'sd588, 32'sd1500, 32'sd877,
32'sd1957, 32'sd1884, 32'sd1756, 32'sd1087, 32'sd1088, 32'sd477,
32'sd119, 32'sd1816, 32'sd1473, 32'sd1906, 32'sd1572, 32'sd1038,
32'sd1151, 32'sd233, 32'sd1690, 32'sd1050, 32'sd1862, 32'sd416,
32'sd1326, 32'sd1181, 32'sd1183, 32'sd886, 32'sd1910, 32'sd1070,
32'sd382, 32'sd1005, 32'sd1662, 32'sd1417, 32'sd680, 32'sd1276,
32'sd671, 32'sd1680, 32'sd954, 32'sd696, 32'sd777, 32'sd604,
32'sd122, 32'sd1496, 32'sd1135, 32'sd1965, 32'sd1406, 32'sd1042,
32'sd1027, 32'sd182, 32'sd484, 32'sd963, 32'sd1439, 32'sd1920,
32'sd581, 32'sd818, 32'sd1943, 32'sd1169, 32'sd1125, 32'sd1592,
32'sd1169, 32'sd375, 32'sd1969, 32'sd719, 32'sd1296, 32'sd1938,
32'sd1909, 32'sd278, 32'sd1582, 32'sd1692, 32'sd772, 32'sd1995,
32'sd857, 32'sd575, 32'sd395, 32'sd1649, 32'sd1969, 32'sd402,
32'sd1750, 32'sd1773, 32'sd459, 32'sd1324, 32'sd1088, 32'sd241,
32'sd850, 32'sd839, 32'sd1540, 32'sd1000, 32'sd1765, 32'sd1016,
32'sd1290, 32'sd965, 32'sd384, 32'sd1233, 32'sd887, 32'sd417,
32'sd1275, 32'sd1429, 32'sd1694, 32'sd1655, 32'sd1284, 32'sd923,
32'sd352, 32'sd1599, 32'sd555, 32'sd147, 32'sd1222, 32'sd383,
32'sd1820, 32'sd1058, 32'sd957, 32'sd1655, 32'sd1130, 32'sd1492,
32'sd1144, 32'sd695, 32'sd1657, 32'sd401, 32'sd637, 32'sd783,
32'sd1435, 32'sd1927, 32'sd1406, 32'sd1178, 32'sd192, 32'sd1945,
32'sd290, 32'sd343, 32'sd1742, 32'sd1126, 32'sd1408, 32'sd266,
32'sd938, 32'sd777, 32'sd245, 32'sd670, 32'sd1801, 32'sd1926,
32'sd1614, 32'sd1647, 32'sd1894, 32'sd1539, 32'sd863, 32'sd600,
32'sd176, 32'sd1398, 32'sd1547, 32'sd885, 32'sd198, 32'sd1940,
32'sd1889, 32'sd302, 32'sd1182, 32'sd182, 32'sd1001, 32'sd1997,
32'sd1335, 32'sd417, 32'sd1655, 32'sd1598, 32'sd1500, 32'sd487,
32'sd803, 32'sd323, 32'sd1025, 32'sd1362, 32'sd440, 32'sd1593,
32'sd1093, 32'sd1765, 32'sd1638, 32'sd1839, 32'sd512, 32'sd311,
32'sd368, 32'sd1281, 32'sd1150, 32'sd1147, 32'sd555, 32'sd444,
32'sd1775, 32'sd234, 32'sd510, 32'sd1130, 32'sd1115, 32'sd971,
32'sd925, 32'sd353, 32'sd226, 32'sd1933, 32'sd1757, 32'sd461,
32'sd1436, 32'sd1771, 32'sd943, 32'sd1274, 32'sd752, 32'sd1752,
32'sd1573, 32'sd340, 32'sd1655, 32'sd1005, 32'sd1760, 32'sd1500,
32'sd1382, 32'sd332, 32'sd988, 32'sd1498, 32'sd1408, 32'sd1959,
32'sd363, 32'sd114, 32'sd1824, 32'sd1840, 32'sd1452, 32'sd1421,
32'sd1969, 32'sd849, 32'sd1020, 32'sd637, 32'sd1811, 32'sd1172,
32'sd842, 32'sd1747, 32'sd829, 32'sd1606, 32'sd1788, 32'sd924,
32'sd1868, 32'sd499, 32'sd981, 32'sd594, 32'sd1239, 32'sd556,
32'sd319, 32'sd1384, 32'sd765, 32'sd765, 32'sd497, 32'sd1619,
32'sd752, 32'sd1898, 32'sd347, 32'sd158, 32'sd904, 32'sd1791,
32'sd1851, 32'sd1662, 32'sd438, 32'sd1770, 32'sd1879, 32'sd336,
32'sd798, 32'sd807, 32'sd1782, 32'sd1302, 32'sd252, 32'sd418,
32'sd1668, 32'sd899, 32'sd1546, 32'sd1113, 32'sd107, 32'sd968,
32'sd199, 32'sd652, 32'sd1555, 32'sd777, 32'sd396, 32'sd1321,
32'sd1827, 32'sd590, 32'sd685, 32'sd315, 32'sd1036, 32'sd1554,
32'sd1703, 32'sd1007, 32'sd163, 32'sd771, 32'sd162, 32'sd693,
32'sd1082, 32'sd1121, 32'sd697, 32'sd1222, 32'sd280, 32'sd708,
32'sd1001, 32'sd1000, 32'sd320, 32'sd513, 32'sd538, 32'sd980,
32'sd398, 32'sd184, 32'sd829, 32'sd1625, 32'sd1467, 32'sd417,
32'sd1731, 32'sd359, 32'sd784, 32'sd1372, 32'sd776, 32'sd870,
32'sd1767, 32'sd785, 32'sd1718, 32'sd1466, 32'sd1033, 32'sd119,
32'sd954, 32'sd1917, 32'sd1237, 32'sd1642, 32'sd965, 32'sd642,
32'sd855, 32'sd499, 32'sd1452, 32'sd550, 32'sd827, 32'sd1496,
32'sd1323, 32'sd620, 32'sd1987, 32'sd1238, 32'sd833, 32'sd855,
32'sd1290, 32'sd1549, 32'sd1678, 32'sd1058, 32'sd1646, 32'sd1847,
32'sd1048, 32'sd356, 32'sd383, 32'sd418, 32'sd191, 32'sd106,
32'sd1100, 32'sd1930, 32'sd1470, 32'sd1167, 32'sd1199, 32'sd1496,
32'sd391, 32'sd601, 32'sd1037, 32'sd583, 32'sd815, 32'sd882,
32'sd711, 32'sd1608, 32'sd1370, 32'sd1620, 32'sd253, 32'sd827,
32'sd328, 32'sd1890, 32'sd1831, 32'sd350, 32'sd1640, 32'sd171,
32'sd859, 32'sd1277, 32'sd1289, 32'sd228, 32'sd1702, 32'sd339,
32'sd865, 32'sd1787, 32'sd1048, 32'sd1372, 32'sd1937, 32'sd1761,
32'sd538, 32'sd1657, 32'sd1963, 32'sd781, 32'sd338, 32'sd1941,
32'sd403, 32'sd1404, 32'sd219, 32'sd936, 32'sd508, 32'sd1742,
32'sd833, 32'sd602, 32'sd714, 32'sd534, 32'sd1636, 32'sd1403,
32'sd872, 32'sd562, 32'sd1808, 32'sd125, 32'sd723, 32'sd112,
32'sd1861, 32'sd708, 32'sd469, 32'sd1558, 32'sd940, 32'sd568,
32'sd125, 32'sd1508, 32'sd475, 32'sd807, 32'sd271, 32'sd617,
32'sd1872, 32'sd885, 32'sd1717, 32'sd1582, 32'sd1289, 32'sd381,
32'sd1707, 32'sd1791, 32'sd1113, 32'sd390, 32'sd629, 32'sd860,
32'sd274, 32'sd1583, 32'sd1192, 32'sd1671, 32'sd1851, 32'sd1377,
32'sd1484, 32'sd171, 32'sd1791, 32'sd1245, 32'sd139, 32'sd1771,
32'sd828, 32'sd1494, 32'sd1197, 32'sd1270, 32'sd1716, 32'sd1686,
32'sd217, 32'sd720, 32'sd505, 32'sd798, 32'sd1158, 32'sd133,
32'sd1103, 32'sd246, 32'sd1072, 32'sd920, 32'sd1671, 32'sd216,
32'sd1054, 32'sd409, 32'sd1002, 32'sd1542, 32'sd411, 32'sd188,
32'sd1767, 32'sd489, 32'sd338, 32'sd565, 32'sd737, 32'sd312,
32'sd1485, 32'sd901, 32'sd1467, 32'sd1466, 32'sd1492, 32'sd571,
32'sd1380, 32'sd683, 32'sd642, 32'sd144, 32'sd1051, 32'sd623,
32'sd1044, 32'sd737, 32'sd1816, 32'sd1403, 32'sd373, 32'sd1893,
32'sd199, 32'sd370, 32'sd1126, 32'sd1708, 32'sd1320, 32'sd1952,
32'sd1026, 32'sd967, 32'sd961, 32'sd1037, 32'sd1006, 32'sd1466,
32'sd334, 32'sd312, 32'sd1925, 32'sd1236, 32'sd1666, 32'sd888,
32'sd1164, 32'sd939, 32'sd390, 32'sd546, 32'sd1579, 32'sd1467,
32'sd1867, 32'sd1546, 32'sd1649, 32'sd1175, 32'sd717, 32'sd101,
32'sd1128, 32'sd565, 32'sd1488, 32'sd1078, 32'sd1395, 32'sd129,
32'sd987, 32'sd628, 32'sd1393, 32'sd1798, 32'sd1608, 32'sd1055,
32'sd525, 32'sd785, 32'sd211, 32'sd660, 32'sd1977, 32'sd1112,
32'sd1954, 32'sd1205, 32'sd1457, 32'sd652, 32'sd852, 32'sd1354,
32'sd689, 32'sd549, 32'sd715, 32'sd1128, 32'sd460, 32'sd248,
32'sd498, 32'sd1028, 32'sd442, 32'sd1073, 32'sd180, 32'sd782,
32'sd135, 32'sd1423, 32'sd1860, 32'sd729, 32'sd1113, 32'sd1828,
32'sd1877, 32'sd984, 32'sd1769, 32'sd141, 32'sd511, 32'sd1493,
32'sd1670, 32'sd1476, 32'sd229, 32'sd293, 32'sd596, 32'sd1130,
32'sd449, 32'sd1391, 32'sd1371, 32'sd375, 32'sd1077, 32'sd1160,
32'sd855, 32'sd1723, 32'sd1486, 32'sd331, 32'sd475, 32'sd115,
32'sd650, 32'sd194, 32'sd232, 32'sd513, 32'sd700, 32'sd1494,
32'sd203, 32'sd932, 32'sd1284, 32'sd185, 32'sd1730, 32'sd829,
32'sd1523, 32'sd182, 32'sd1581, 32'sd701, 32'sd429, 32'sd830,
32'sd1189, 32'sd1415, 32'sd1840, 32'sd1995, 32'sd1369, 32'sd120,
32'sd908, 32'sd308, 32'sd798, 32'sd1034, 32'sd965, 32'sd1693,
32'sd353, 32'sd1704, 32'sd194, 32'sd507, 32'sd346, 32'sd1244,
32'sd735, 32'sd1405, 32'sd1793, 32'sd1840, 32'sd1750, 32'sd1035,
32'sd1931, 32'sd414, 32'sd1107, 32'sd1018, 32'sd1987, 32'sd1956,
32'sd1224, 32'sd914, 32'sd708, 32'sd1432, 32'sd1283, 32'sd1440,
32'sd1823, 32'sd851, 32'sd500, 32'sd630, 32'sd123, 32'sd760,
32'sd530, 32'sd1218, 32'sd300, 32'sd876, 32'sd949, 32'sd1857,
32'sd1683, 32'sd1892, 32'sd1026, 32'sd1386, 32'sd1391, 32'sd1742,
32'sd1145, 32'sd1631, 32'sd570, 32'sd1090, 32'sd573, 32'sd105,
32'sd701, 32'sd1708, 32'sd1422, 32'sd1489, 32'sd1063, 32'sd1513,
32'sd1107, 32'sd1250, 32'sd1662, 32'sd885, 32'sd427, 32'sd195,
32'sd1146, 32'sd257, 32'sd1077, 32'sd807, 32'sd230, 32'sd1512,
32'sd785, 32'sd299, 32'sd551, 32'sd506, 32'sd110, 32'sd1683,
32'sd365, 32'sd851, 32'sd1077, 32'sd1919, 32'sd1058, 32'sd1067,
32'sd1962, 32'sd1049, 32'sd1681, 32'sd1250, 32'sd1058, 32'sd246,
32'sd473, 32'sd304, 32'sd745, 32'sd1567, 32'sd149, 32'sd832,
32'sd844, 32'sd327, 32'sd1985, 32'sd401, 32'sd1738, 32'sd145,
32'sd884, 32'sd1743, 32'sd814, 32'sd865, 32'sd1451, 32'sd1664,
32'sd245, 32'sd1402, 32'sd444, 32'sd273, 32'sd278, 32'sd889,
32'sd1623, 32'sd1848, 32'sd1007, 32'sd1865, 32'sd1857, 32'sd1602,
32'sd1996, 32'sd1762, 32'sd1588, 32'sd1011, 32'sd1835, 32'sd1566,
32'sd557, 32'sd471, 32'sd912, 32'sd812, 32'sd1088, 32'sd1020,
32'sd725, 32'sd1824, 32'sd1552, 32'sd1440, 32'sd1771, 32'sd1611,
32'sd191, 32'sd318, 32'sd1023, 32'sd1028, 32'sd539, 32'sd850,
32'sd570, 32'sd584, 32'sd527, 32'sd1124, 32'sd1766, 32'sd1915,
32'sd465, 32'sd929, 32'sd1289, 32'sd1231, 32'sd1823, 32'sd1489,
32'sd384, 32'sd167, 32'sd1471, 32'sd1628, 32'sd1590, 32'sd1462,
32'sd1068, 32'sd243, 32'sd1355, 32'sd1329, 32'sd1157, 32'sd1587,
32'sd569, 32'sd1140, 32'sd1787, 32'sd1050, 32'sd1190, 32'sd336,
32'sd1661, 32'sd1759, 32'sd367, 32'sd1391, 32'sd650, 32'sd1324,
32'sd1628, 32'sd1127, 32'sd273, 32'sd221, 32'sd1824, 32'sd1788,
32'sd1849, 32'sd289, 32'sd1518, 32'sd1521, 32'sd1791, 32'sd552,
32'sd921, 32'sd786, 32'sd624, 32'sd1789, 32'sd1085, 32'sd210,
32'sd988, 32'sd794, 32'sd878, 32'sd903, 32'sd768, 32'sd1857,
32'sd664, 32'sd1205, 32'sd309, 32'sd232, 32'sd374, 32'sd1952,
32'sd249, 32'sd1376, 32'sd637, 32'sd1619, 32'sd1557, 32'sd1824,
32'sd1924, 32'sd1245, 32'sd847, 32'sd1131, 32'sd876, 32'sd1431,
32'sd297, 32'sd1083, 32'sd844, 32'sd1767, 32'sd1005, 32'sd1995,
32'sd925, 32'sd772, 32'sd193, 32'sd805, 32'sd119, 32'sd1000,
32'sd782, 32'sd420, 32'sd1857, 32'sd1234, 32'sd1768, 32'sd1744,
32'sd1722, 32'sd875, 32'sd1633, 32'sd1644, 32'sd1889, 32'sd1997,
32'sd1329, 32'sd1723, 32'sd189, 32'sd125, 32'sd1295, 32'sd790,
32'sd300, 32'sd1697, 32'sd1610, 32'sd221, 32'sd1961, 32'sd478,
32'sd1199, 32'sd1833, 32'sd542, 32'sd218, 32'sd195, 32'sd1587,
32'sd1701, 32'sd1656, 32'sd1914, 32'sd421, 32'sd1094, 32'sd912,
32'sd1441, 32'sd1861, 32'sd931, 32'sd152, 32'sd1437, 32'sd766,
32'sd663, 32'sd1989, 32'sd1730, 32'sd936, 32'sd1614, 32'sd711,
32'sd1360, 32'sd1621, 32'sd506, 32'sd424, 32'sd1775, 32'sd412,
32'sd774, 32'sd1813, 32'sd1426, 32'sd581, 32'sd1268, 32'sd1469,
32'sd1689, 32'sd574, 32'sd1680, 32'sd1529, 32'sd1841, 32'sd1522,
32'sd1833, 32'sd1706, 32'sd1050, 32'sd1038, 32'sd1239, 32'sd635,
32'sd694, 32'sd1704, 32'sd1486, 32'sd128, 32'sd1563, 32'sd846,
32'sd1631, 32'sd1137, 32'sd1475, 32'sd1398, 32'sd137, 32'sd835,
32'sd1650, 32'sd1511, 32'sd970, 32'sd363, 32'sd288, 32'sd807,
32'sd1078, 32'sd986, 32'sd427, 32'sd1019, 32'sd1480, 32'sd1165,
32'sd1013, 32'sd1143, 32'sd427, 32'sd444, 32'sd557, 32'sd1399,
32'sd1401, 32'sd826, 32'sd1462, 32'sd133, 32'sd103, 32'sd568,
32'sd661, 32'sd1009, 32'sd711, 32'sd425, 32'sd1180, 32'sd591,
32'sd1562, 32'sd1260, 32'sd821, 32'sd220, 32'sd643, 32'sd157,
32'sd1125, 32'sd277, 32'sd1187, 32'sd591, 32'sd1453, 32'sd757,
32'sd289, 32'sd1527, 32'sd1093, 32'sd204, 32'sd1107, 32'sd109,
32'sd1363, 32'sd449, 32'sd1912, 32'sd1647, 32'sd1503, 32'sd1801,
32'sd1687, 32'sd1829, 32'sd695, 32'sd1424, 32'sd1270, 32'sd637,
32'sd1716, 32'sd425, 32'sd420, 32'sd961, 32'sd1300, 32'sd1966,
32'sd1710, 32'sd697, 32'sd313, 32'sd154, 32'sd1388, 32'sd175,
32'sd1070, 32'sd735, 32'sd1877, 32'sd403, 32'sd1047, 32'sd202,
32'sd868, 32'sd579, 32'sd1518, 32'sd927, 32'sd1482, 32'sd1194,
32'sd1142, 32'sd1314, 32'sd860, 32'sd608, 32'sd1406, 32'sd1252,
32'sd618, 32'sd237, 32'sd768, 32'sd1190, 32'sd1257, 32'sd280,
32'sd795, 32'sd1430, 32'sd337, 32'sd732, 32'sd1317, 32'sd964,
32'sd497, 32'sd1267, 32'sd334, 32'sd283, 32'sd1670, 32'sd1923,
32'sd224, 32'sd1332, 32'sd1874, 32'sd489, 32'sd621, 32'sd432,
32'sd643, 32'sd1538, 32'sd946, 32'sd187, 32'sd1972, 32'sd918,
32'sd651, 32'sd1518, 32'sd760, 32'sd1291, 32'sd1941, 32'sd1210,
32'sd937, 32'sd1220, 32'sd352, 32'sd1440, 32'sd109, 32'sd724,
32'sd726, 32'sd254, 32'sd448, 32'sd1524, 32'sd173, 32'sd1461,
32'sd1117, 32'sd1768, 32'sd1749, 32'sd1497, 32'sd1458, 32'sd1597,
32'sd1697, 32'sd324, 32'sd1802, 32'sd791, 32'sd1649, 32'sd1887,
32'sd689, 32'sd621, 32'sd1326, 32'sd1373, 32'sd588, 32'sd1289,
32'sd430, 32'sd1542, 32'sd259, 32'sd1228, 32'sd794, 32'sd1666,
32'sd799, 32'sd1606, 32'sd1590, 32'sd358, 32'sd1617, 32'sd1833,
32'sd1790, 32'sd1087, 32'sd225, 32'sd1239, 32'sd901, 32'sd1814,
32'sd1273, 32'sd1598, 32'sd1659, 32'sd945, 32'sd1979, 32'sd973,
32'sd855, 32'sd1557, 32'sd1817, 32'sd1643, 32'sd1860, 32'sd762,
32'sd499, 32'sd233, 32'sd1406, 32'sd1403, 32'sd996, 32'sd174,
32'sd989, 32'sd889, 32'sd741, 32'sd1908, 32'sd540, 32'sd571,
32'sd903, 32'sd1445, 32'sd695, 32'sd176, 32'sd1263, 32'sd1317,
32'sd1184, 32'sd1994, 32'sd940, 32'sd352, 32'sd269, 32'sd820,
32'sd1295, 32'sd1639, 32'sd306, 32'sd1294, 32'sd1749, 32'sd1381,
32'sd1784, 32'sd1562, 32'sd935, 32'sd634, 32'sd1504, 32'sd1272,
32'sd1718, 32'sd1428, 32'sd1313, 32'sd1777, 32'sd1138, 32'sd1874,
32'sd1570, 32'sd369, 32'sd1772, 32'sd432, 32'sd1509, 32'sd989,
32'sd1078, 32'sd1390, 32'sd1686, 32'sd1405, 32'sd1538, 32'sd1923,
32'sd101, 32'sd1862, 32'sd1069, 32'sd1969, 32'sd439, 32'sd1213,
32'sd349, 32'sd1213, 32'sd1322, 32'sd1392, 32'sd1438, 32'sd280,
32'sd1522, 32'sd1648, 32'sd536, 32'sd536, 32'sd1484, 32'sd146,
32'sd1591, 32'sd1011, 32'sd1326, 32'sd1830, 32'sd263, 32'sd157,
32'sd1418, 32'sd1650, 32'sd1783, 32'sd934, 32'sd1388, 32'sd1062,
32'sd666, 32'sd143, 32'sd948, 32'sd774, 32'sd944, 32'sd1161,
32'sd328, 32'sd941, 32'sd608, 32'sd871, 32'sd424, 32'sd1713,
32'sd169, 32'sd1705, 32'sd1089, 32'sd1085, 32'sd1361, 32'sd852,
32'sd1546, 32'sd1361, 32'sd678, 32'sd850, 32'sd795, 32'sd761,
32'sd374, 32'sd205, 32'sd1066, 32'sd119, 32'sd1256, 32'sd1383,
32'sd712, 32'sd930, 32'sd1600, 32'sd873, 32'sd778, 32'sd1670,
32'sd1802, 32'sd1343, 32'sd1736, 32'sd889, 32'sd1926, 32'sd606,
32'sd530, 32'sd391, 32'sd344, 32'sd1822, 32'sd847, 32'sd462,
32'sd1374, 32'sd1107, 32'sd321, 32'sd1935, 32'sd1953, 32'sd293,
32'sd555, 32'sd1929, 32'sd1567, 32'sd850, 32'sd1553, 32'sd1777,
32'sd1687, 32'sd261, 32'sd682, 32'sd406, 32'sd862, 32'sd1664,
32'sd522, 32'sd263, 32'sd239, 32'sd1306, 32'sd664, 32'sd1107,
32'sd504, 32'sd1199, 32'sd1135, 32'sd664, 32'sd175, 32'sd834,
32'sd552, 32'sd726, 32'sd1619, 32'sd1565, 32'sd957, 32'sd651,
32'sd1641, 32'sd1327, 32'sd665, 32'sd1501, 32'sd1200, 32'sd990,
32'sd546, 32'sd1166, 32'sd906, 32'sd224, 32'sd1951, 32'sd248,
32'sd196, 32'sd451, 32'sd1365, 32'sd439, 32'sd822, 32'sd1502,
32'sd1183, 32'sd656, 32'sd275, 32'sd390, 32'sd235, 32'sd1435,
32'sd1667, 32'sd886, 32'sd626, 32'sd1243, 32'sd1101, 32'sd524,
32'sd1836, 32'sd1787, 32'sd1410, 32'sd684, 32'sd1829, 32'sd352,
32'sd765, 32'sd1578, 32'sd765, 32'sd921, 32'sd512, 32'sd711,
32'sd1535, 32'sd487, 32'sd1519, 32'sd1163, 32'sd1533, 32'sd1876,
32'sd1194, 32'sd1227, 32'sd1157, 32'sd924, 32'sd1349, 32'sd505,
32'sd549, 32'sd675, 32'sd1604, 32'sd500, 32'sd243, 32'sd771,
32'sd100, 32'sd288, 32'sd1588, 32'sd1290, 32'sd1895, 32'sd1233,
32'sd1549, 32'sd873, 32'sd601, 32'sd239, 32'sd1195, 32'sd1253,
32'sd1033, 32'sd994, 32'sd1747, 32'sd346, 32'sd1690, 32'sd510,
32'sd1083, 32'sd1649, 32'sd1208, 32'sd1427, 32'sd1039, 32'sd1689,
32'sd998, 32'sd909, 32'sd1879, 32'sd127, 32'sd286, 32'sd1293,
32'sd432, 32'sd736, 32'sd1297, 32'sd1055, 32'sd1374, 32'sd1079,
32'sd1068, 32'sd313, 32'sd1695, 32'sd1987, 32'sd1945, 32'sd638,
32'sd1026, 32'sd1789, 32'sd1060, 32'sd305, 32'sd166, 32'sd849,
32'sd747, 32'sd586, 32'sd1368, 32'sd1259, 32'sd1558, 32'sd1427,
32'sd1673, 32'sd1424, 32'sd1644, 32'sd1207, 32'sd427, 32'sd1901,
32'sd298, 32'sd1518, 32'sd416, 32'sd898, 32'sd366, 32'sd1369,
32'sd1453, 32'sd140, 32'sd437, 32'sd290, 32'sd1740, 32'sd1161,
32'sd120, 32'sd1081, 32'sd1062, 32'sd1108, 32'sd321, 32'sd1296,
32'sd875, 32'sd311, 32'sd1706, 32'sd136, 32'sd640, 32'sd1273,
32'sd1665, 32'sd129, 32'sd1906, 32'sd310, 32'sd306, 32'sd1635,
32'sd1628, 32'sd1267, 32'sd599, 32'sd1478, 32'sd1987, 32'sd350,
32'sd470, 32'sd1980, 32'sd1530, 32'sd179, 32'sd1275, 32'sd1378,
32'sd106, 32'sd1417, 32'sd1298, 32'sd1665, 32'sd381, 32'sd915,
32'sd1575, 32'sd465, 32'sd1509, 32'sd620, 32'sd826, 32'sd1138,
32'sd932, 32'sd1451, 32'sd1113, 32'sd1562, 32'sd1937, 32'sd428,
32'sd1758, 32'sd1807, 32'sd1857, 32'sd1582, 32'sd1733, 32'sd1214,
32'sd1804, 32'sd1922, 32'sd1202, 32'sd1159, 32'sd193, 32'sd1149,
32'sd307, 32'sd1367, 32'sd1875, 32'sd1344, 32'sd410, 32'sd1501,
32'sd1009, 32'sd786, 32'sd635, 32'sd943, 32'sd119, 32'sd1322,
32'sd843, 32'sd960, 32'sd854, 32'sd614, 32'sd158, 32'sd1674,
32'sd1773, 32'sd1192, 32'sd500, 32'sd1817, 32'sd114, 32'sd626,
32'sd1648, 32'sd372, 32'sd641, 32'sd1584, 32'sd1686, 32'sd1002,
32'sd1459, 32'sd655, 32'sd1193, 32'sd393, 32'sd726, 32'sd917,
32'sd1187, 32'sd496, 32'sd1377, 32'sd1608, 32'sd1596, 32'sd720,
32'sd869, 32'sd803, 32'sd1680, 32'sd1695, 32'sd1983, 32'sd1186,
32'sd1485, 32'sd779, 32'sd1631, 32'sd854, 32'sd1020, 32'sd1674,
32'sd582, 32'sd939, 32'sd737, 32'sd1290, 32'sd1236, 32'sd1719,
32'sd736, 32'sd626, 32'sd1788, 32'sd1494, 32'sd835, 32'sd1690,
32'sd797, 32'sd1561, 32'sd1674, 32'sd601, 32'sd1912, 32'sd1692,
32'sd1939, 32'sd853, 32'sd1193, 32'sd1355, 32'sd562, 32'sd693,
32'sd1302, 32'sd1250, 32'sd1014, 32'sd167, 32'sd1015, 32'sd860,
32'sd1744, 32'sd707, 32'sd1164, 32'sd1707, 32'sd1854, 32'sd1642,
32'sd110, 32'sd1979, 32'sd527, 32'sd1751, 32'sd300, 32'sd1790,
32'sd1603, 32'sd1279, 32'sd629, 32'sd1251, 32'sd869, 32'sd1272,
32'sd1657, 32'sd449, 32'sd1135, 32'sd1237, 32'sd1565, 32'sd902,
32'sd1337, 32'sd251, 32'sd427, 32'sd673, 32'sd1566, 32'sd1372,
32'sd1850, 32'sd620, 32'sd913, 32'sd1672, 32'sd844, 32'sd958,
32'sd1762, 32'sd717, 32'sd881, 32'sd1754, 32'sd829, 32'sd900,
32'sd443, 32'sd1433, 32'sd1876, 32'sd1614, 32'sd960, 32'sd1755,
32'sd1803, 32'sd1432, 32'sd409, 32'sd1840, 32'sd839, 32'sd1207,
32'sd361, 32'sd837, 32'sd1839, 32'sd1714, 32'sd1187, 32'sd288,
32'sd1206, 32'sd540, 32'sd359, 32'sd412, 32'sd1403, 32'sd1265,
32'sd1040, 32'sd670, 32'sd1569, 32'sd140, 32'sd1350, 32'sd1761,
32'sd1153, 32'sd1165, 32'sd1933, 32'sd1499, 32'sd574, 32'sd1796,
32'sd1000, 32'sd901, 32'sd538, 32'sd197, 32'sd185, 32'sd1234,
32'sd1827, 32'sd1981, 32'sd1558, 32'sd971, 32'sd358, 32'sd1363,
32'sd284, 32'sd1083, 32'sd1545, 32'sd1664, 32'sd839, 32'sd341,
32'sd1414, 32'sd115, 32'sd1746, 32'sd663, 32'sd1422, 32'sd850,
32'sd821, 32'sd1195, 32'sd1622, 32'sd1213, 32'sd1126, 32'sd1727,
32'sd207, 32'sd1712, 32'sd672, 32'sd1115, 32'sd1880, 32'sd608,
32'sd210, 32'sd1310, 32'sd945, 32'sd1680, 32'sd1246, 32'sd1149,
32'sd1544, 32'sd887, 32'sd102, 32'sd1475, 32'sd1637, 32'sd335,
32'sd896, 32'sd1353, 32'sd540, 32'sd765, 32'sd521, 32'sd124,
32'sd1213, 32'sd1611, 32'sd1892, 32'sd1295, 32'sd1641, 32'sd1619,
32'sd1981, 32'sd846, 32'sd1914, 32'sd1209, 32'sd1217, 32'sd910,
32'sd1310, 32'sd1830, 32'sd788, 32'sd1624, 32'sd610, 32'sd847,
32'sd1690, 32'sd528, 32'sd1027, 32'sd1707, 32'sd1541, 32'sd690,
32'sd1381, 32'sd699, 32'sd1846, 32'sd1184, 32'sd476, 32'sd1456,
32'sd1949, 32'sd1051, 32'sd1246, 32'sd1839, 32'sd1496, 32'sd1066,
32'sd1058, 32'sd545, 32'sd457, 32'sd1226, 32'sd1263, 32'sd1699,
32'sd1047, 32'sd1030, 32'sd1709, 32'sd1531, 32'sd1862, 32'sd1994,
32'sd189, 32'sd879, 32'sd746, 32'sd1525, 32'sd1243, 32'sd468,
32'sd961, 32'sd1071, 32'sd1620, 32'sd214, 32'sd1510, 32'sd593,
32'sd621, 32'sd453, 32'sd160, 32'sd790, 32'sd1275, 32'sd1812,
32'sd558, 32'sd1313, 32'sd515, 32'sd1708, 32'sd1233, 32'sd677,
32'sd1401, 32'sd1638, 32'sd1747, 32'sd735, 32'sd654, 32'sd1824,
32'sd1191, 32'sd642, 32'sd1424, 32'sd1025, 32'sd1255, 32'sd1287,
32'sd1721, 32'sd1867, 32'sd750, 32'sd855, 32'sd689, 32'sd1390,
32'sd406, 32'sd1279, 32'sd557, 32'sd196, 32'sd263, 32'sd962,
32'sd1811, 32'sd1248, 32'sd1159, 32'sd337, 32'sd291, 32'sd701,
32'sd700, 32'sd649, 32'sd366, 32'sd1948, 32'sd1239, 32'sd781,
32'sd625, 32'sd1712, 32'sd446, 32'sd341, 32'sd1126, 32'sd1434,
32'sd552, 32'sd855, 32'sd745, 32'sd383, 32'sd1156, 32'sd598,
32'sd309, 32'sd231, 32'sd1527, 32'sd752, 32'sd1969, 32'sd1470,
32'sd570, 32'sd556, 32'sd1201, 32'sd902, 32'sd1016, 32'sd479,
32'sd858, 32'sd1556, 32'sd316, 32'sd923, 32'sd122, 32'sd773,
32'sd513, 32'sd1287, 32'sd1757, 32'sd842, 32'sd718, 32'sd830,
32'sd196, 32'sd653, 32'sd711, 32'sd134, 32'sd1486, 32'sd1290,
32'sd614, 32'sd1249, 32'sd1586, 32'sd1867, 32'sd989, 32'sd1260,
32'sd1175, 32'sd1049, 32'sd1689, 32'sd1225, 32'sd1813, 32'sd788,
32'sd929, 32'sd1497, 32'sd529, 32'sd143, 32'sd1724, 32'sd972,
32'sd1273, 32'sd1682, 32'sd1141, 32'sd1556, 32'sd1491, 32'sd1359,
32'sd247, 32'sd1518, 32'sd642, 32'sd616, 32'sd648, 32'sd743,
32'sd635, 32'sd758, 32'sd945, 32'sd279, 32'sd1774, 32'sd1074,
32'sd1281, 32'sd670, 32'sd306, 32'sd838, 32'sd1485, 32'sd1907,
32'sd1132, 32'sd1238, 32'sd792, 32'sd292, 32'sd1612, 32'sd1361,
32'sd629, 32'sd815, 32'sd653, 32'sd237, 32'sd105, 32'sd472,
32'sd1589, 32'sd695, 32'sd475, 32'sd458, 32'sd1712, 32'sd667,
32'sd246, 32'sd722, 32'sd1118, 32'sd494, 32'sd355, 32'sd110,
32'sd1247, 32'sd649, 32'sd974, 32'sd1961, 32'sd253, 32'sd507,
32'sd500, 32'sd1786, 32'sd1222, 32'sd411, 32'sd1209, 32'sd1567,
32'sd808, 32'sd1600, 32'sd1028, 32'sd1528, 32'sd1822, 32'sd1467,
32'sd947, 32'sd1341, 32'sd1551, 32'sd685, 32'sd1336, 32'sd808,
32'sd1906, 32'sd1712, 32'sd230, 32'sd1585, 32'sd1448, 32'sd1434,
32'sd133, 32'sd920, 32'sd332, 32'sd1115, 32'sd1578, 32'sd837,
32'sd1925, 32'sd1186, 32'sd170, 32'sd1031, 32'sd1590, 32'sd1957,
32'sd659, 32'sd220, 32'sd630, 32'sd1848, 32'sd379, 32'sd1886,
32'sd1635, 32'sd1804, 32'sd140, 32'sd1598, 32'sd1102, 32'sd1332,
32'sd1341, 32'sd1698, 32'sd1079, 32'sd414, 32'sd950, 32'sd777,
32'sd1339, 32'sd1194, 32'sd1128, 32'sd1571, 32'sd1715, 32'sd734,
32'sd152, 32'sd168, 32'sd119, 32'sd1083, 32'sd812, 32'sd1811,
32'sd1049, 32'sd1462, 32'sd1593, 32'sd1361, 32'sd1840, 32'sd178,
32'sd695, 32'sd1012, 32'sd752, 32'sd127, 32'sd533, 32'sd904,
32'sd843, 32'sd1494, 32'sd1155, 32'sd1857, 32'sd1682, 32'sd530,
32'sd443, 32'sd190, 32'sd1624, 32'sd1682, 32'sd1733, 32'sd1153,
32'sd1933, 32'sd1060, 32'sd860, 32'sd572, 32'sd222, 32'sd456,
32'sd1877, 32'sd1623, 32'sd349, 32'sd1649, 32'sd1235, 32'sd1130,
32'sd1326, 32'sd649, 32'sd663, 32'sd1670, 32'sd1937, 32'sd104,
32'sd814, 32'sd1348, 32'sd752, 32'sd431, 32'sd974, 32'sd1872,
32'sd742, 32'sd996, 32'sd1302, 32'sd120, 32'sd1701, 32'sd601,
32'sd993, 32'sd550, 32'sd1714, 32'sd810, 32'sd1310, 32'sd857,
32'sd360, 32'sd252, 32'sd563, 32'sd439, 32'sd473, 32'sd280,
32'sd1276, 32'sd244, 32'sd690, 32'sd761, 32'sd1519, 32'sd1629,
32'sd467, 32'sd451, 32'sd113, 32'sd180, 32'sd1590, 32'sd1822,
32'sd1937, 32'sd722, 32'sd141, 32'sd1660, 32'sd775, 32'sd1117,
32'sd1091, 32'sd1928, 32'sd158, 32'sd1572, 32'sd479, 32'sd1864,
32'sd1380, 32'sd1050, 32'sd1595, 32'sd1557, 32'sd1440, 32'sd423,
32'sd1332, 32'sd641, 32'sd1148, 32'sd1922, 32'sd130, 32'sd347,
32'sd636, 32'sd768, 32'sd1712, 32'sd501, 32'sd963, 32'sd386,
32'sd192, 32'sd1023, 32'sd719, 32'sd345, 32'sd1569, 32'sd1935,
32'sd386, 32'sd2000, 32'sd1602, 32'sd1099, 32'sd1287, 32'sd1663,
32'sd1940, 32'sd1561, 32'sd1477, 32'sd267, 32'sd1885, 32'sd1852,
32'sd719, 32'sd1589, 32'sd1801, 32'sd870, 32'sd176, 32'sd1486,
32'sd710, 32'sd771, 32'sd1547, 32'sd741, 32'sd1283, 32'sd809,
32'sd683, 32'sd1128, 32'sd1693, 32'sd871, 32'sd387, 32'sd721,
32'sd1560, 32'sd749, 32'sd1949, 32'sd248, 32'sd1926, 32'sd546,
32'sd1948, 32'sd135, 32'sd1125, 32'sd1494, 32'sd1494, 32'sd781,
32'sd1460, 32'sd635, 32'sd1334, 32'sd1594, 32'sd693, 32'sd170,
32'sd1330, 32'sd1877, 32'sd294, 32'sd1079, 32'sd748, 32'sd113,
32'sd1872, 32'sd316, 32'sd1903, 32'sd895, 32'sd556, 32'sd1275,
32'sd758, 32'sd663, 32'sd1826, 32'sd1604, 32'sd1202, 32'sd1753,
32'sd1638, 32'sd1048, 32'sd1498, 32'sd895, 32'sd1470, 32'sd761,
32'sd1378, 32'sd1165, 32'sd1250, 32'sd744, 32'sd757, 32'sd871,
32'sd1834, 32'sd833, 32'sd1403, 32'sd733, 32'sd753, 32'sd1965,
32'sd1318, 32'sd1069, 32'sd1851, 32'sd642, 32'sd155, 32'sd1321,
32'sd1573, 32'sd604, 32'sd1174, 32'sd1783, 32'sd1879, 32'sd1525,
32'sd1346, 32'sd1094, 32'sd1230, 32'sd1937, 32'sd170, 32'sd1134,
32'sd140, 32'sd1725, 32'sd169, 32'sd1036, 32'sd1973, 32'sd1833,
32'sd1546, 32'sd629, 32'sd1831, 32'sd1236, 32'sd862, 32'sd492,
32'sd1501, 32'sd1751, 32'sd1089, 32'sd1362, 32'sd2000, 32'sd1372,
32'sd1864, 32'sd1746, 32'sd1169, 32'sd1262, 32'sd529, 32'sd556,
32'sd1025, 32'sd278, 32'sd867, 32'sd1232, 32'sd1065, 32'sd1386,
32'sd1338, 32'sd659, 32'sd366, 32'sd962, 32'sd1233, 32'sd453,
32'sd786, 32'sd1392, 32'sd1702, 32'sd845, 32'sd760, 32'sd1176,
32'sd406, 32'sd1101, 32'sd129, 32'sd705, 32'sd124, 32'sd1561,
32'sd1376, 32'sd1682, 32'sd588, 32'sd1323, 32'sd1724, 32'sd1418,
32'sd989, 32'sd444, 32'sd1786, 32'sd1081, 32'sd820, 32'sd682,
32'sd419, 32'sd940, 32'sd144, 32'sd1765, 32'sd998, 32'sd466,
32'sd799, 32'sd1471, 32'sd498, 32'sd1227, 32'sd1616, 32'sd871,
32'sd1617, 32'sd1404, 32'sd1461, 32'sd627, 32'sd1583, 32'sd223,
32'sd1919, 32'sd319, 32'sd406, 32'sd753, 32'sd1540, 32'sd1206,
32'sd1437, 32'sd1441, 32'sd1846, 32'sd364, 32'sd1040, 32'sd1708,
32'sd937, 32'sd371, 32'sd581, 32'sd1665, 32'sd1777, 32'sd1862,
32'sd550, 32'sd1978, 32'sd850, 32'sd1819, 32'sd1888, 32'sd289,
32'sd827, 32'sd531, 32'sd809, 32'sd1279, 32'sd597, 32'sd516,
32'sd1322, 32'sd1332, 32'sd851, 32'sd1830, 32'sd1259, 32'sd190,
32'sd211, 32'sd1552, 32'sd574, 32'sd1722, 32'sd712, 32'sd977,
32'sd1841, 32'sd349, 32'sd766, 32'sd1610, 32'sd1427, 32'sd638,
32'sd1224, 32'sd437, 32'sd569, 32'sd1946, 32'sd1719, 32'sd1540,
32'sd1233, 32'sd1000, 32'sd1962, 32'sd1561, 32'sd1474, 32'sd104,
32'sd1258, 32'sd498, 32'sd1421, 32'sd573, 32'sd1450, 32'sd1319,
32'sd350, 32'sd291, 32'sd894, 32'sd1400, 32'sd1125, 32'sd1635,
32'sd1772, 32'sd1553, 32'sd423, 32'sd1827, 32'sd628, 32'sd434,
32'sd542, 32'sd1200, 32'sd1516, 32'sd169, 32'sd167, 32'sd134,
32'sd1470, 32'sd1851, 32'sd1809, 32'sd1253, 32'sd668, 32'sd1017,
32'sd1216, 32'sd1906, 32'sd1394, 32'sd651, 32'sd172, 32'sd1515,
32'sd879, 32'sd1033, 32'sd312, 32'sd874, 32'sd296, 32'sd805,
32'sd1089, 32'sd954, 32'sd885, 32'sd1084, 32'sd1295, 32'sd1879,
32'sd335, 32'sd604, 32'sd1586, 32'sd1035, 32'sd1718, 32'sd1229,
32'sd1281, 32'sd631, 32'sd509, 32'sd1702, 32'sd624, 32'sd1999,
32'sd994, 32'sd1564, 32'sd707, 32'sd1525, 32'sd1427, 32'sd1079,
32'sd1735, 32'sd759, 32'sd1228, 32'sd1094, 32'sd1993, 32'sd588,
32'sd724, 32'sd521, 32'sd1215, 32'sd1559, 32'sd799, 32'sd950,
32'sd615, 32'sd1544, 32'sd1725, 32'sd1322, 32'sd554, 32'sd1962,
32'sd906, 32'sd905, 32'sd1486, 32'sd719, 32'sd1823, 32'sd307,
32'sd2000, 32'sd1022, 32'sd904, 32'sd1329, 32'sd1333, 32'sd291,
32'sd1032, 32'sd489, 32'sd1001, 32'sd447, 32'sd918, 32'sd809,
32'sd841, 32'sd799, 32'sd808, 32'sd689, 32'sd1507, 32'sd1236,
32'sd1572, 32'sd557, 32'sd613, 32'sd1897, 32'sd742, 32'sd1661,
32'sd468, 32'sd1928, 32'sd358, 32'sd587, 32'sd793, 32'sd591,
32'sd1438, 32'sd1520, 32'sd1768, 32'sd674, 32'sd1125, 32'sd1722,
32'sd982, 32'sd1334, 32'sd655, 32'sd1038, 32'sd223, 32'sd1392,
32'sd218, 32'sd932, 32'sd116, 32'sd1730, 32'sd429, 32'sd1251,
32'sd995, 32'sd637, 32'sd1976, 32'sd1275, 32'sd1804, 32'sd1928,
32'sd1759, 32'sd1341, 32'sd1781, 32'sd816, 32'sd1939, 32'sd442,
32'sd1662, 32'sd535, 32'sd1242, 32'sd630, 32'sd1478, 32'sd1425,
32'sd1954, 32'sd1515, 32'sd1986, 32'sd1813, 32'sd1241, 32'sd457,
32'sd1349, 32'sd396, 32'sd209, 32'sd379, 32'sd1262, 32'sd1000,
32'sd1898, 32'sd1947, 32'sd1803, 32'sd1223, 32'sd1103, 32'sd158,
32'sd568, 32'sd203, 32'sd1204, 32'sd1797, 32'sd391, 32'sd706,
32'sd284, 32'sd1764, 32'sd1180, 32'sd1496, 32'sd1736, 32'sd378,
32'sd1682, 32'sd1710, 32'sd697, 32'sd1025, 32'sd1835, 32'sd1767,
32'sd399, 32'sd1366, 32'sd1756, 32'sd672, 32'sd909, 32'sd214,
32'sd126, 32'sd1900, 32'sd859, 32'sd238, 32'sd719, 32'sd1225,
32'sd354, 32'sd1700, 32'sd1570, 32'sd144, 32'sd756, 32'sd1618,
32'sd835, 32'sd1299, 32'sd335, 32'sd1198, 32'sd721, 32'sd536,
32'sd1981, 32'sd1302, 32'sd1040, 32'sd199, 32'sd274, 32'sd1612,
32'sd1760, 32'sd1098, 32'sd620, 32'sd1855, 32'sd1180, 32'sd116,
32'sd1769, 32'sd290, 32'sd251, 32'sd1037, 32'sd787, 32'sd1466,
32'sd1634, 32'sd1077, 32'sd984, 32'sd1556, 32'sd226, 32'sd396,
32'sd751, 32'sd1623, 32'sd1604, 32'sd1931, 32'sd1108, 32'sd1752,
32'sd250, 32'sd1345, 32'sd1443, 32'sd995, 32'sd153, 32'sd1954,
32'sd1105, 32'sd292, 32'sd978, 32'sd438, 32'sd592, 32'sd303,
32'sd1284, 32'sd1239, 32'sd518, 32'sd1397, 32'sd1826, 32'sd443,
32'sd627, 32'sd743, 32'sd1039, 32'sd1257, 32'sd219, 32'sd1799,
32'sd529, 32'sd1314, 32'sd797, 32'sd1126, 32'sd1700, 32'sd686,
32'sd1644, 32'sd1477, 32'sd403, 32'sd361, 32'sd1992, 32'sd1135,
32'sd1735, 32'sd562, 32'sd1039, 32'sd490, 32'sd765, 32'sd1924,
32'sd367, 32'sd1034, 32'sd1267, 32'sd666, 32'sd416, 32'sd1932,
32'sd258, 32'sd304, 32'sd773, 32'sd1216, 32'sd1055, 32'sd1250,
32'sd1192, 32'sd1261, 32'sd546, 32'sd906, 32'sd287, 32'sd775,
32'sd1315, 32'sd1424, 32'sd288, 32'sd1722, 32'sd1659, 32'sd188,
32'sd497, 32'sd1022, 32'sd1235, 32'sd812, 32'sd1037, 32'sd528,
32'sd506, 32'sd1303, 32'sd1481, 32'sd1338, 32'sd1336, 32'sd767,
32'sd1480, 32'sd1480, 32'sd1417, 32'sd805, 32'sd911, 32'sd920,
32'sd425, 32'sd1664, 32'sd227, 32'sd1176, 32'sd1216, 32'sd1058,
32'sd1877, 32'sd269, 32'sd1075, 32'sd866, 32'sd1544, 32'sd1930,
32'sd278, 32'sd1754, 32'sd1889, 32'sd687, 32'sd1768, 32'sd1719,
32'sd228, 32'sd1907, 32'sd1292, 32'sd875, 32'sd951, 32'sd546,
32'sd475, 32'sd1952, 32'sd1134, 32'sd1029, 32'sd252, 32'sd1384,
32'sd325, 32'sd403, 32'sd247, 32'sd668, 32'sd756, 32'sd552,
32'sd720, 32'sd413, 32'sd1486, 32'sd334, 32'sd1071, 32'sd765,
32'sd942, 32'sd1648, 32'sd1062, 32'sd396, 32'sd628, 32'sd790,
32'sd558, 32'sd1640, 32'sd812, 32'sd1536, 32'sd1976, 32'sd661,
32'sd1049, 32'sd1733, 32'sd655, 32'sd1094, 32'sd134, 32'sd1081,
32'sd992, 32'sd1618, 32'sd530, 32'sd495, 32'sd113, 32'sd709,
32'sd1555, 32'sd1988, 32'sd1519, 32'sd1919, 32'sd705, 32'sd868,
32'sd214, 32'sd1785, 32'sd297, 32'sd1658, 32'sd1140, 32'sd717,
32'sd1250, 32'sd861, 32'sd1030, 32'sd1537, 32'sd1063, 32'sd210,
32'sd1673, 32'sd487, 32'sd1482, 32'sd482, 32'sd171, 32'sd1597,
32'sd213, 32'sd702, 32'sd1443, 32'sd1357, 32'sd1963, 32'sd625,
32'sd1636, 32'sd1021, 32'sd170, 32'sd289, 32'sd1082, 32'sd1411,
32'sd234, 32'sd1024, 32'sd1243, 32'sd149, 32'sd1689, 32'sd1805,
32'sd152, 32'sd1563, 32'sd244, 32'sd1946, 32'sd800, 32'sd1744,
32'sd980, 32'sd401, 32'sd1606, 32'sd1108, 32'sd726, 32'sd783,
32'sd924, 32'sd1446, 32'sd696, 32'sd1620, 32'sd1057, 32'sd474,
32'sd678, 32'sd282, 32'sd1483, 32'sd657, 32'sd1893, 32'sd728,
32'sd1266, 32'sd582, 32'sd1144, 32'sd976, 32'sd844, 32'sd1278,
32'sd932, 32'sd1269, 32'sd509, 32'sd1521, 32'sd881, 32'sd1754,
32'sd1570, 32'sd978, 32'sd1181, 32'sd282, 32'sd210, 32'sd289,
32'sd154, 32'sd535, 32'sd1859, 32'sd1076, 32'sd1103, 32'sd1856,
32'sd1809, 32'sd1899, 32'sd587, 32'sd305, 32'sd1978, 32'sd980,
32'sd1907, 32'sd805, 32'sd1274, 32'sd440, 32'sd928, 32'sd1690,
32'sd1860, 32'sd1936, 32'sd886, 32'sd804, 32'sd1941, 32'sd731,
32'sd230, 32'sd130, 32'sd1931, 32'sd1561, 32'sd1645, 32'sd323,
32'sd670, 32'sd790, 32'sd406, 32'sd1769, 32'sd421, 32'sd1189,
32'sd347, 32'sd695, 32'sd1815, 32'sd236, 32'sd1877, 32'sd556,
32'sd1858, 32'sd1604, 32'sd500, 32'sd1137, 32'sd440, 32'sd1760,
32'sd1962, 32'sd687, 32'sd1689, 32'sd832, 32'sd1817, 32'sd1659,
32'sd1848, 32'sd1764, 32'sd1651, 32'sd1857, 32'sd161, 32'sd235,
32'sd1538, 32'sd1912, 32'sd463, 32'sd941, 32'sd242, 32'sd1636,
32'sd908, 32'sd1574, 32'sd514, 32'sd1926, 32'sd1359, 32'sd1538,
32'sd799, 32'sd1123, 32'sd1901, 32'sd1708, 32'sd1420, 32'sd1765,
32'sd1376, 32'sd741, 32'sd507, 32'sd1588, 32'sd1975, 32'sd215,
32'sd1958, 32'sd258, 32'sd442, 32'sd185, 32'sd1206, 32'sd1226,
32'sd477, 32'sd1135, 32'sd146, 32'sd1258, 32'sd1993, 32'sd222,
32'sd283, 32'sd487, 32'sd1989, 32'sd987, 32'sd1338, 32'sd1004,
32'sd1838, 32'sd1720, 32'sd1992, 32'sd225, 32'sd1215, 32'sd419,
32'sd1010, 32'sd1018, 32'sd832, 32'sd393, 32'sd199, 32'sd1545,
32'sd982, 32'sd170, 32'sd1803, 32'sd647, 32'sd1859, 32'sd1512,
32'sd1103, 32'sd521, 32'sd1997, 32'sd742, 32'sd928, 32'sd333,
32'sd356, 32'sd722, 32'sd764, 32'sd813, 32'sd206, 32'sd1373,
32'sd111, 32'sd351, 32'sd126, 32'sd623, 32'sd880, 32'sd1421,
32'sd1755, 32'sd1348, 32'sd579, 32'sd1610, 32'sd725, 32'sd1800,
32'sd1198, 32'sd1929, 32'sd614, 32'sd1099, 32'sd360, 32'sd1799,
32'sd1011, 32'sd496, 32'sd169, 32'sd1613, 32'sd337, 32'sd844,
32'sd1921, 32'sd571, 32'sd611, 32'sd1656, 32'sd157, 32'sd1449,
32'sd1836, 32'sd307, 32'sd1601, 32'sd1047, 32'sd1219, 32'sd448,
32'sd503, 32'sd1621, 32'sd1413, 32'sd1919, 32'sd244, 32'sd1311,
32'sd1402, 32'sd694, 32'sd1804, 32'sd1101, 32'sd207, 32'sd1477,
32'sd716, 32'sd1321, 32'sd628, 32'sd1661, 32'sd925, 32'sd868,
32'sd857, 32'sd673, 32'sd874, 32'sd1321, 32'sd951, 32'sd1357,
32'sd814, 32'sd1973, 32'sd476, 32'sd1104, 32'sd559, 32'sd386,
32'sd669, 32'sd100, 32'sd796, 32'sd1308, 32'sd1022, 32'sd439,
32'sd694, 32'sd181, 32'sd878, 32'sd947, 32'sd834, 32'sd587,
32'sd1876, 32'sd366, 32'sd500, 32'sd205, 32'sd1444, 32'sd1036,
32'sd657, 32'sd1719, 32'sd635, 32'sd779, 32'sd698, 32'sd514,
32'sd239, 32'sd1679, 32'sd119, 32'sd485, 32'sd154, 32'sd1810,
32'sd193, 32'sd1238, 32'sd997, 32'sd756, 32'sd1568, 32'sd1182,
32'sd278, 32'sd1328, 32'sd744, 32'sd232, 32'sd1316, 32'sd666,
32'sd756, 32'sd176, 32'sd1580, 32'sd1580, 32'sd1665, 32'sd1219,
32'sd1089, 32'sd1116, 32'sd572, 32'sd1164, 32'sd1372, 32'sd639,
32'sd1240, 32'sd1989, 32'sd923, 32'sd791, 32'sd1458, 32'sd1883,
32'sd1582, 32'sd1419, 32'sd1443, 32'sd1257, 32'sd754, 32'sd1079,
32'sd349, 32'sd741, 32'sd652, 32'sd1326, 32'sd1977, 32'sd877,
32'sd1125, 32'sd793, 32'sd1298, 32'sd203, 32'sd246, 32'sd961,
32'sd1971, 32'sd1714, 32'sd1435, 32'sd602, 32'sd1756, 32'sd1920,
32'sd1274, 32'sd1642, 32'sd786, 32'sd156, 32'sd1898, 32'sd1651,
32'sd1073, 32'sd1091, 32'sd243, 32'sd858, 32'sd685, 32'sd1648,
32'sd1995, 32'sd1254, 32'sd103, 32'sd1936, 32'sd1528, 32'sd1585,
32'sd725, 32'sd1603, 32'sd1914, 32'sd1180, 32'sd748, 32'sd621,
32'sd1561, 32'sd759, 32'sd1076, 32'sd1967, 32'sd306, 32'sd1775,
32'sd1656, 32'sd1360, 32'sd193, 32'sd1520, 32'sd517, 32'sd926,
32'sd330, 32'sd152, 32'sd748, 32'sd745, 32'sd1042, 32'sd276,
32'sd1005, 32'sd1713, 32'sd577, 32'sd1589, 32'sd1729, 32'sd1237,
32'sd770, 32'sd1249, 32'sd310, 32'sd1629, 32'sd1158, 32'sd1775,
32'sd1558, 32'sd807, 32'sd1795, 32'sd1056, 32'sd1722, 32'sd1283,
32'sd1347, 32'sd1767, 32'sd1457, 32'sd992, 32'sd297, 32'sd1980,
32'sd390, 32'sd1704, 32'sd891, 32'sd965, 32'sd185, 32'sd1862,
32'sd1630, 32'sd285, 32'sd1697, 32'sd1413, 32'sd400, 32'sd1905,
32'sd1721, 32'sd1999, 32'sd968, 32'sd370, 32'sd1961, 32'sd1437,
32'sd1659, 32'sd1902, 32'sd1396, 32'sd167, 32'sd1648, 32'sd1072,
32'sd883, 32'sd831, 32'sd221, 32'sd776, 32'sd1170, 32'sd667,
32'sd291, 32'sd528, 32'sd1502, 32'sd1074, 32'sd1147, 32'sd1887,
32'sd1473, 32'sd1042, 32'sd1076, 32'sd906, 32'sd810, 32'sd1964,
32'sd1336, 32'sd1409, 32'sd1714, 32'sd1531, 32'sd752, 32'sd1922,
32'sd671, 32'sd406, 32'sd1020, 32'sd276, 32'sd1129, 32'sd1724,
32'sd1388, 32'sd1167, 32'sd1389, 32'sd1351, 32'sd1854, 32'sd1155,
32'sd647, 32'sd1231, 32'sd1032, 32'sd1776, 32'sd1996, 32'sd1298,
32'sd1134, 32'sd1440, 32'sd291, 32'sd911, 32'sd375, 32'sd1251,
32'sd794, 32'sd754, 32'sd1985, 32'sd842, 32'sd732, 32'sd1751,
32'sd365, 32'sd969, 32'sd1086, 32'sd1397, 32'sd725, 32'sd196,
32'sd1480, 32'sd130, 32'sd688, 32'sd802, 32'sd632, 32'sd108,
32'sd1958, 32'sd1332, 32'sd766, 32'sd509, 32'sd288, 32'sd1020,
32'sd934, 32'sd1995, 32'sd523, 32'sd1711, 32'sd1684, 32'sd881,
32'sd1789, 32'sd226, 32'sd428, 32'sd764, 32'sd1483, 32'sd603,
32'sd1351, 32'sd1005, 32'sd1995, 32'sd1411, 32'sd920, 32'sd144,
32'sd1632, 32'sd222, 32'sd389, 32'sd446, 32'sd1310, 32'sd267,
32'sd708, 32'sd1848, 32'sd1519, 32'sd1105, 32'sd481, 32'sd967,
32'sd131, 32'sd650, 32'sd1547, 32'sd317, 32'sd1786, 32'sd1306,
32'sd613, 32'sd1614, 32'sd473, 32'sd1399, 32'sd944, 32'sd1776,
32'sd1878, 32'sd115, 32'sd1070, 32'sd1949, 32'sd826, 32'sd724,
32'sd817, 32'sd808, 32'sd186, 32'sd1756, 32'sd557, 32'sd1571,
32'sd693, 32'sd1210, 32'sd617, 32'sd1192, 32'sd758, 32'sd930,
32'sd664, 32'sd1644, 32'sd1079, 32'sd770, 32'sd1904, 32'sd1371,
32'sd1809, 32'sd878, 32'sd445, 32'sd604, 32'sd587, 32'sd1904,
32'sd1810, 32'sd1474, 32'sd193, 32'sd985, 32'sd285, 32'sd1665,
32'sd1763, 32'sd634, 32'sd1776, 32'sd395, 32'sd1533, 32'sd1172,
32'sd903, 32'sd799, 32'sd927, 32'sd1614, 32'sd772, 32'sd1684,
32'sd1472, 32'sd802, 32'sd1121, 32'sd884, 32'sd885, 32'sd199,
32'sd423, 32'sd190, 32'sd1943, 32'sd702, 32'sd851, 32'sd1572,
32'sd906, 32'sd1071, 32'sd1769, 32'sd938, 32'sd513, 32'sd1531,
32'sd1322, 32'sd1416, 32'sd118, 32'sd1944, 32'sd130, 32'sd1798,
32'sd965, 32'sd1508, 32'sd1546, 32'sd196, 32'sd257, 32'sd949,
32'sd378, 32'sd1569, 32'sd1968, 32'sd925, 32'sd799, 32'sd1938,
32'sd766, 32'sd1902, 32'sd216, 32'sd543, 32'sd1118, 32'sd667,
32'sd1951, 32'sd950, 32'sd792, 32'sd1684, 32'sd220, 32'sd1403,
32'sd256, 32'sd1928, 32'sd1594, 32'sd874, 32'sd1507, 32'sd1131,
32'sd1671, 32'sd909, 32'sd1532, 32'sd1783, 32'sd1076, 32'sd1568,
32'sd1175, 32'sd445, 32'sd431, 32'sd1079, 32'sd315, 32'sd1356,
32'sd1163, 32'sd1759, 32'sd326, 32'sd818, 32'sd397, 32'sd988,
32'sd1521, 32'sd440, 32'sd1964, 32'sd314, 32'sd1549, 32'sd1800,
32'sd545, 32'sd383, 32'sd1206, 32'sd833, 32'sd1481, 32'sd939,
32'sd1154, 32'sd914, 32'sd1664, 32'sd314, 32'sd101, 32'sd1720,
32'sd1746, 32'sd439, 32'sd127, 32'sd118, 32'sd1093, 32'sd816,
32'sd507, 32'sd558, 32'sd809, 32'sd1204, 32'sd341, 32'sd292,
32'sd1442, 32'sd525, 32'sd1452, 32'sd406, 32'sd1968, 32'sd1114,
32'sd248, 32'sd687, 32'sd1733, 32'sd901, 32'sd243, 32'sd1839,
32'sd319, 32'sd500, 32'sd398, 32'sd832, 32'sd1954, 32'sd1804,
32'sd1848, 32'sd198, 32'sd1322, 32'sd1149, 32'sd922, 32'sd1841,
32'sd1763, 32'sd673, 32'sd1898, 32'sd1164, 32'sd1977, 32'sd1210,
32'sd1931, 32'sd654, 32'sd1372, 32'sd1540, 32'sd803, 32'sd873,
32'sd1739, 32'sd401, 32'sd1662, 32'sd1539, 32'sd1576, 32'sd1200,
32'sd1398, 32'sd1904, 32'sd850, 32'sd983, 32'sd1532, 32'sd315,
32'sd1452, 32'sd959, 32'sd1113, 32'sd262, 32'sd385, 32'sd519,
32'sd132, 32'sd1783, 32'sd1471, 32'sd1022, 32'sd1037, 32'sd1384,
32'sd1788, 32'sd109, 32'sd912, 32'sd1845, 32'sd961, 32'sd977,
32'sd1784, 32'sd1987, 32'sd1542, 32'sd498, 32'sd1621, 32'sd1087,
32'sd282, 32'sd910, 32'sd1223, 32'sd1950, 32'sd574, 32'sd1895,
32'sd651, 32'sd538, 32'sd1713, 32'sd1949, 32'sd1429, 32'sd606,
32'sd1126, 32'sd166, 32'sd1740, 32'sd182, 32'sd1109, 32'sd1539,
32'sd1339, 32'sd1153, 32'sd1696, 32'sd806, 32'sd1264, 32'sd793,
32'sd1640, 32'sd1403, 32'sd1096, 32'sd222, 32'sd1087, 32'sd1231,
32'sd1303, 32'sd572, 32'sd1254, 32'sd1780, 32'sd1324, 32'sd285,
32'sd631, 32'sd548, 32'sd1173, 32'sd861, 32'sd246, 32'sd615,
32'sd1127, 32'sd1702, 32'sd839, 32'sd1253, 32'sd770, 32'sd595,
32'sd1782, 32'sd1588, 32'sd115, 32'sd1533, 32'sd702, 32'sd1361,
32'sd128, 32'sd1015, 32'sd1377, 32'sd305, 32'sd1922, 32'sd1787,
32'sd1711, 32'sd1216, 32'sd1711, 32'sd622, 32'sd471, 32'sd1606,
32'sd1989, 32'sd1251, 32'sd1662, 32'sd1275, 32'sd875, 32'sd368,
32'sd1185, 32'sd1041, 32'sd256, 32'sd692, 32'sd663, 32'sd688,
32'sd252, 32'sd1969, 32'sd1498, 32'sd225, 32'sd1735, 32'sd208,
32'sd1977, 32'sd634, 32'sd1617, 32'sd1864, 32'sd1415, 32'sd594,
32'sd1662, 32'sd512, 32'sd110, 32'sd1202, 32'sd361, 32'sd1595,
32'sd1488, 32'sd1290, 32'sd1912, 32'sd1151, 32'sd1801, 32'sd960,
32'sd217, 32'sd752, 32'sd1062, 32'sd1496, 32'sd1932, 32'sd1522,
32'sd502, 32'sd383, 32'sd1191, 32'sd1607, 32'sd1276, 32'sd1968,
32'sd1943, 32'sd327, 32'sd1537, 32'sd1492, 32'sd1847, 32'sd1497,
32'sd288, 32'sd789, 32'sd1381, 32'sd348, 32'sd1481, 32'sd1773,
32'sd1181, 32'sd1351, 32'sd1597, 32'sd975, 32'sd1814, 32'sd591,
32'sd223, 32'sd1369, 32'sd1115, 32'sd1006, 32'sd1623, 32'sd577,
32'sd377, 32'sd1623, 32'sd1932, 32'sd242, 32'sd981, 32'sd573,
32'sd1905, 32'sd733, 32'sd1974, 32'sd812, 32'sd113, 32'sd458,
32'sd1645, 32'sd617, 32'sd630, 32'sd756, 32'sd1390, 32'sd1233,
32'sd1989, 32'sd236, 32'sd588, 32'sd1471, 32'sd1201, 32'sd964,
32'sd884, 32'sd848, 32'sd1391, 32'sd1728, 32'sd1110, 32'sd1300,
32'sd1720, 32'sd140, 32'sd1610, 32'sd1447, 32'sd296, 32'sd2000,
32'sd1789, 32'sd1704, 32'sd444, 32'sd976, 32'sd1408, 32'sd1318,
32'sd1746, 32'sd1589, 32'sd1976, 32'sd539, 32'sd510, 32'sd584,
32'sd165, 32'sd1941, 32'sd1002, 32'sd1231, 32'sd1848, 32'sd1201,
32'sd1870, 32'sd650, 32'sd1798, 32'sd1769, 32'sd494, 32'sd130,
32'sd1191, 32'sd782, 32'sd856, 32'sd1938, 32'sd674, 32'sd976,
32'sd1575, 32'sd1836, 32'sd1463, 32'sd961, 32'sd216, 32'sd1288,
32'sd238, 32'sd277, 32'sd1646, 32'sd228, 32'sd195, 32'sd140,
32'sd1691, 32'sd1768, 32'sd1893, 32'sd1832, 32'sd653, 32'sd462,
32'sd1522, 32'sd1578, 32'sd368, 32'sd1389, 32'sd1230, 32'sd606,
32'sd1688, 32'sd1797, 32'sd1594, 32'sd688, 32'sd941, 32'sd722,
32'sd513, 32'sd139, 32'sd909, 32'sd560, 32'sd1670, 32'sd1551,
32'sd799, 32'sd366, 32'sd796, 32'sd1856, 32'sd1911, 32'sd1717,
32'sd987, 32'sd1235, 32'sd100, 32'sd122, 32'sd128, 32'sd1415,
32'sd1084, 32'sd734, 32'sd1313, 32'sd1943, 32'sd424, 32'sd498,
32'sd1702, 32'sd537, 32'sd965, 32'sd1502, 32'sd501, 32'sd1924,
32'sd1623, 32'sd701, 32'sd877, 32'sd1674, 32'sd967, 32'sd1405,
32'sd1835, 32'sd624, 32'sd1868, 32'sd198, 32'sd635, 32'sd774,
32'sd501, 32'sd757, 32'sd1298, 32'sd143, 32'sd141, 32'sd996,
32'sd709, 32'sd906, 32'sd629, 32'sd1058, 32'sd1257, 32'sd1256,
32'sd1203, 32'sd1335, 32'sd1424, 32'sd970, 32'sd494, 32'sd803,
32'sd762, 32'sd1281, 32'sd1507, 32'sd391, 32'sd1376, 32'sd492,
32'sd316, 32'sd1904, 32'sd1285, 32'sd1459, 32'sd1500, 32'sd1311,
32'sd1124, 32'sd1199, 32'sd1413, 32'sd497, 32'sd272, 32'sd1887,
32'sd869, 32'sd450, 32'sd1245, 32'sd230, 32'sd1658, 32'sd812,
32'sd1862, 32'sd1177, 32'sd372, 32'sd987, 32'sd502, 32'sd758,
32'sd1423, 32'sd514, 32'sd874, 32'sd1762, 32'sd1700, 32'sd1900,
32'sd1695, 32'sd189, 32'sd237, 32'sd629, 32'sd702, 32'sd1022,
32'sd280, 32'sd986, 32'sd1915, 32'sd914, 32'sd1819, 32'sd1625,
32'sd1796, 32'sd1480, 32'sd697, 32'sd421, 32'sd589, 32'sd1323,
32'sd447, 32'sd252, 32'sd390, 32'sd730, 32'sd1713, 32'sd1463,
32'sd1005, 32'sd1526, 32'sd1203, 32'sd1421, 32'sd1732, 32'sd987,
32'sd1370, 32'sd873, 32'sd352, 32'sd823, 32'sd120, 32'sd1204,
32'sd1922, 32'sd1654, 32'sd1459, 32'sd1225, 32'sd956, 32'sd209,
32'sd1070, 32'sd1917, 32'sd1286, 32'sd1158, 32'sd474, 32'sd362,
32'sd574, 32'sd749, 32'sd1734, 32'sd1409, 32'sd204, 32'sd1358,
32'sd110, 32'sd1932, 32'sd1568, 32'sd1602, 32'sd418, 32'sd924,
32'sd603, 32'sd1706, 32'sd222, 32'sd1993, 32'sd1990, 32'sd852,
32'sd1586, 32'sd1732, 32'sd1456, 32'sd591, 32'sd1300, 32'sd1675,
32'sd205, 32'sd1704, 32'sd1861, 32'sd248, 32'sd1960, 32'sd116,
32'sd552, 32'sd325, 32'sd1833, 32'sd785, 32'sd1155, 32'sd195,
32'sd1186, 32'sd402, 32'sd225, 32'sd162, 32'sd1177, 32'sd100,
32'sd1437, 32'sd632, 32'sd1289, 32'sd1237, 32'sd1765, 32'sd179,
32'sd629, 32'sd1888, 32'sd1640, 32'sd1099, 32'sd518, 32'sd1328,
32'sd770, 32'sd1395, 32'sd204, 32'sd618, 32'sd692, 32'sd1819,
32'sd1811, 32'sd1206, 32'sd1691, 32'sd1344, 32'sd1223, 32'sd1124,
32'sd1733, 32'sd716, 32'sd1796, 32'sd329, 32'sd1309, 32'sd1095,
32'sd1190, 32'sd1406, 32'sd1033, 32'sd1771, 32'sd109, 32'sd1703,
32'sd185, 32'sd1298, 32'sd1609, 32'sd588, 32'sd1608, 32'sd348,
32'sd791, 32'sd350, 32'sd466, 32'sd517, 32'sd1798, 32'sd376,
32'sd1555, 32'sd613, 32'sd793, 32'sd566, 32'sd375, 32'sd304,
32'sd1149, 32'sd1518, 32'sd1533, 32'sd1967, 32'sd1944, 32'sd518,
32'sd1881, 32'sd555, 32'sd194, 32'sd961, 32'sd1384, 32'sd817,
32'sd185, 32'sd1810, 32'sd1458, 32'sd1172, 32'sd436, 32'sd169,
32'sd587, 32'sd996, 32'sd1111, 32'sd541, 32'sd797, 32'sd1949,
32'sd177, 32'sd822, 32'sd771, 32'sd692, 32'sd1260, 32'sd1387,
32'sd111, 32'sd1191, 32'sd1810, 32'sd1920, 32'sd1062, 32'sd552,
32'sd108, 32'sd213, 32'sd1471, 32'sd1782, 32'sd1910, 32'sd943,
32'sd1203, 32'sd297, 32'sd1043, 32'sd1317, 32'sd1386, 32'sd367,
32'sd1435, 32'sd741, 32'sd1627, 32'sd707, 32'sd117, 32'sd1119,
32'sd1847, 32'sd1448, 32'sd1392, 32'sd795, 32'sd1113, 32'sd1025,
32'sd557, 32'sd1825, 32'sd133, 32'sd1357, 32'sd497, 32'sd276,
32'sd1335, 32'sd1459, 32'sd834, 32'sd1289, 32'sd965, 32'sd1466,
32'sd779, 32'sd1733, 32'sd1414, 32'sd134, 32'sd1199, 32'sd1398,
32'sd233, 32'sd998, 32'sd1672, 32'sd267, 32'sd1069, 32'sd954,
32'sd915, 32'sd1631, 32'sd1354, 32'sd634, 32'sd213, 32'sd875,
32'sd566, 32'sd993, 32'sd1743, 32'sd192, 32'sd355, 32'sd363,
32'sd1077, 32'sd1972, 32'sd126, 32'sd309, 32'sd186, 32'sd863,
32'sd1746, 32'sd643, 32'sd1865, 32'sd937, 32'sd1326, 32'sd1654,
32'sd1959, 32'sd1208, 32'sd935, 32'sd887, 32'sd1275, 32'sd1337,
32'sd1800, 32'sd1220, 32'sd482, 32'sd604, 32'sd703, 32'sd1756,
32'sd545, 32'sd209, 32'sd1807, 32'sd1794, 32'sd902, 32'sd1704,
32'sd1948, 32'sd1104, 32'sd286, 32'sd1218, 32'sd109, 32'sd709,
32'sd682, 32'sd113, 32'sd617, 32'sd1602, 32'sd819, 32'sd1758,
32'sd829, 32'sd1117, 32'sd1512, 32'sd1255, 32'sd554, 32'sd1938,
32'sd1398, 32'sd1736, 32'sd805, 32'sd949, 32'sd542, 32'sd479,
32'sd747, 32'sd1913, 32'sd946, 32'sd1869, 32'sd1509, 32'sd1054,
32'sd1467, 32'sd742, 32'sd1561, 32'sd1416, 32'sd969, 32'sd1711,
32'sd1770, 32'sd333, 32'sd786, 32'sd174, 32'sd913, 32'sd517,
32'sd409, 32'sd1729, 32'sd357, 32'sd832, 32'sd926, 32'sd638,
32'sd761, 32'sd1313, 32'sd1949, 32'sd1312, 32'sd1291, 32'sd488,
32'sd1222, 32'sd795, 32'sd902, 32'sd397, 32'sd1012, 32'sd744,
32'sd1621, 32'sd1416, 32'sd714, 32'sd113, 32'sd1349, 32'sd896,
32'sd1527, 32'sd620, 32'sd1256, 32'sd736, 32'sd761, 32'sd1447,
32'sd184, 32'sd972, 32'sd199, 32'sd871, 32'sd1709, 32'sd1991,
32'sd505, 32'sd1528, 32'sd1204, 32'sd1331, 32'sd223, 32'sd544,
32'sd1891, 32'sd1875, 32'sd1225, 32'sd1250, 32'sd245, 32'sd1384,
32'sd123, 32'sd1889, 32'sd1779, 32'sd630, 32'sd967, 32'sd920,
32'sd1068, 32'sd641, 32'sd124, 32'sd915, 32'sd716, 32'sd1215,
32'sd819, 32'sd589, 32'sd611, 32'sd614, 32'sd644, 32'sd1984,
32'sd317, 32'sd1139, 32'sd439, 32'sd1363, 32'sd1170, 32'sd872,
32'sd1435, 32'sd1009, 32'sd1622, 32'sd1673, 32'sd1008, 32'sd1593,
32'sd507, 32'sd216, 32'sd1792, 32'sd338, 32'sd533, 32'sd222,
32'sd1340, 32'sd869, 32'sd778, 32'sd1434, 32'sd680, 32'sd1592,
32'sd1170, 32'sd291, 32'sd598, 32'sd975, 32'sd1054, 32'sd678,
32'sd1710, 32'sd1710, 32'sd1599, 32'sd896, 32'sd673, 32'sd1960,
32'sd1705, 32'sd1602, 32'sd1692, 32'sd315, 32'sd385, 32'sd634,
32'sd1454, 32'sd1547, 32'sd1241, 32'sd1800, 32'sd1562, 32'sd1363,
32'sd1962, 32'sd349, 32'sd521, 32'sd1920, 32'sd1122, 32'sd1704,
32'sd1120, 32'sd512, 32'sd342, 32'sd184, 32'sd1458, 32'sd1286,
32'sd205, 32'sd167, 32'sd1190, 32'sd747, 32'sd431, 32'sd1928,
32'sd216, 32'sd473, 32'sd637, 32'sd1828, 32'sd590, 32'sd1604,
32'sd1854, 32'sd1304, 32'sd1188, 32'sd1436, 32'sd1310, 32'sd130,
32'sd1717, 32'sd1559, 32'sd1882, 32'sd472, 32'sd1742, 32'sd204,
32'sd740, 32'sd1455, 32'sd985, 32'sd1926, 32'sd327, 32'sd556,
32'sd296, 32'sd1963, 32'sd1212, 32'sd428, 32'sd1883, 32'sd505,
32'sd191, 32'sd1456, 32'sd1675, 32'sd911, 32'sd604, 32'sd1415,
32'sd1258, 32'sd857, 32'sd1483, 32'sd1588, 32'sd1086, 32'sd1070,
32'sd1764, 32'sd1932, 32'sd1343, 32'sd1266, 32'sd1042, 32'sd588,
32'sd1226, 32'sd1142, 32'sd830, 32'sd474, 32'sd711, 32'sd357,
32'sd321, 32'sd1658, 32'sd1023, 32'sd439, 32'sd1658, 32'sd1431,
32'sd742, 32'sd1629, 32'sd1280, 32'sd1696, 32'sd434, 32'sd360,
32'sd1469, 32'sd588, 32'sd1104, 32'sd1934, 32'sd696, 32'sd1655,
32'sd219, 32'sd1861, 32'sd1857, 32'sd694, 32'sd780, 32'sd1740,
32'sd1393, 32'sd636, 32'sd1319, 32'sd919, 32'sd1012, 32'sd1942,
32'sd519, 32'sd1456, 32'sd1542, 32'sd1917, 32'sd1908, 32'sd237,
32'sd561, 32'sd801, 32'sd1358, 32'sd1391, 32'sd718, 32'sd795,
32'sd408, 32'sd282, 32'sd300, 32'sd1043, 32'sd136, 32'sd1282,
32'sd600, 32'sd779, 32'sd278, 32'sd1919, 32'sd1291, 32'sd192,
32'sd1347, 32'sd455, 32'sd1587, 32'sd211, 32'sd227, 32'sd482,
32'sd205, 32'sd905, 32'sd1087, 32'sd399, 32'sd172, 32'sd1551,
32'sd1283, 32'sd354, 32'sd1489, 32'sd150, 32'sd284, 32'sd1888,
32'sd703, 32'sd1808, 32'sd1967, 32'sd1241, 32'sd1681, 32'sd1955,
32'sd1269, 32'sd619, 32'sd1039, 32'sd278, 32'sd237, 32'sd278,
32'sd1057, 32'sd1308, 32'sd799, 32'sd1977, 32'sd937, 32'sd162,
32'sd627, 32'sd1621, 32'sd1109, 32'sd355, 32'sd353, 32'sd1215,
32'sd687, 32'sd1554, 32'sd661, 32'sd278, 32'sd400, 32'sd1636,
32'sd1154, 32'sd1359, 32'sd1764, 32'sd317, 32'sd1881, 32'sd398,
32'sd104, 32'sd551, 32'sd1610, 32'sd1496, 32'sd721, 32'sd260,
32'sd1330, 32'sd534, 32'sd163, 32'sd989, 32'sd1226, 32'sd460,
32'sd1731, 32'sd370, 32'sd936, 32'sd346, 32'sd677, 32'sd427,
32'sd1857, 32'sd910, 32'sd712, 32'sd939, 32'sd1333, 32'sd1942,
32'sd1417, 32'sd424, 32'sd1440, 32'sd1072, 32'sd1876, 32'sd861,
32'sd519, 32'sd206, 32'sd1861, 32'sd1670, 32'sd283, 32'sd847,
32'sd236, 32'sd1800, 32'sd314, 32'sd401, 32'sd821, 32'sd1557,
32'sd283, 32'sd1754, 32'sd1974, 32'sd1688, 32'sd580, 32'sd1589,
32'sd746, 32'sd756, 32'sd1734, 32'sd1945, 32'sd644, 32'sd960,
32'sd349, 32'sd1682, 32'sd1936, 32'sd1414, 32'sd524, 32'sd1552,
32'sd1321, 32'sd522, 32'sd1665, 32'sd112, 32'sd929, 32'sd1814,
32'sd278, 32'sd1010, 32'sd749, 32'sd859, 32'sd535, 32'sd549,
32'sd1148, 32'sd753, 32'sd1916, 32'sd1344, 32'sd715, 32'sd903,
32'sd891, 32'sd966, 32'sd1581, 32'sd1164, 32'sd567, 32'sd139,
32'sd1414, 32'sd1257, 32'sd411, 32'sd1466, 32'sd1847, 32'sd1566,
32'sd1668, 32'sd673, 32'sd715, 32'sd127, 32'sd1301, 32'sd674,
32'sd349, 32'sd769, 32'sd1309, 32'sd359, 32'sd1398, 32'sd436,
32'sd1194, 32'sd427, 32'sd1514, 32'sd708, 32'sd556, 32'sd1848,
32'sd1445, 32'sd1498, 32'sd1882, 32'sd1933, 32'sd878, 32'sd1175,
32'sd547, 32'sd1074, 32'sd988, 32'sd1177, 32'sd920, 32'sd416,
32'sd1422, 32'sd1648, 32'sd589, 32'sd431, 32'sd760, 32'sd1284,
32'sd413, 32'sd1764, 32'sd1776, 32'sd1101, 32'sd1667, 32'sd377,
32'sd748, 32'sd1984, 32'sd1196, 32'sd1230, 32'sd235, 32'sd618,
32'sd480, 32'sd717, 32'sd1102, 32'sd486, 32'sd896, 32'sd1919,
32'sd1094, 32'sd789, 32'sd1487, 32'sd1930, 32'sd582, 32'sd1330,
32'sd1137, 32'sd454, 32'sd624, 32'sd1717, 32'sd746, 32'sd1836,
32'sd1488, 32'sd234, 32'sd1485, 32'sd1956, 32'sd1321, 32'sd1078,
32'sd1297, 32'sd561, 32'sd112, 32'sd604, 32'sd418, 32'sd1582,
32'sd176, 32'sd1499, 32'sd1570, 32'sd1662, 32'sd1591, 32'sd247,
32'sd1020, 32'sd1149, 32'sd408, 32'sd1470, 32'sd1297, 32'sd1210,
32'sd1234, 32'sd612, 32'sd434, 32'sd1941, 32'sd263, 32'sd159,
32'sd1111, 32'sd484, 32'sd941, 32'sd1591, 32'sd1991, 32'sd1900,
32'sd396, 32'sd449, 32'sd1174, 32'sd331, 32'sd290, 32'sd1772,
32'sd1508, 32'sd333, 32'sd230, 32'sd169, 32'sd517, 32'sd1645,
32'sd892, 32'sd1223, 32'sd558, 32'sd753, 32'sd1235, 32'sd550,
32'sd1067, 32'sd1707, 32'sd452, 32'sd498, 32'sd1929, 32'sd989,
32'sd356, 32'sd291, 32'sd395, 32'sd1625, 32'sd1475, 32'sd711,
32'sd1452, 32'sd252, 32'sd681, 32'sd1487, 32'sd1484, 32'sd1168,
32'sd762, 32'sd1482, 32'sd381, 32'sd868, 32'sd1599, 32'sd1272,
32'sd581, 32'sd1296, 32'sd540, 32'sd676, 32'sd1232, 32'sd268,
32'sd1865, 32'sd1628, 32'sd114, 32'sd1633, 32'sd1307, 32'sd312,
32'sd1572, 32'sd612, 32'sd1265, 32'sd523, 32'sd605, 32'sd1026,
32'sd1495, 32'sd1384, 32'sd1625, 32'sd220, 32'sd1521, 32'sd1486,
32'sd1288, 32'sd242, 32'sd1850, 32'sd140, 32'sd1774, 32'sd1565,
32'sd1248, 32'sd1578, 32'sd1410, 32'sd1122, 32'sd1047, 32'sd130,
32'sd1064, 32'sd1731, 32'sd589, 32'sd753, 32'sd335, 32'sd497,
32'sd1775, 32'sd652, 32'sd912, 32'sd310, 32'sd928, 32'sd735,
32'sd1537, 32'sd586, 32'sd250, 32'sd1201, 32'sd325, 32'sd1084,
32'sd1490, 32'sd1949, 32'sd1086, 32'sd1196, 32'sd1493, 32'sd486,
32'sd689, 32'sd989, 32'sd1888, 32'sd750, 32'sd189, 32'sd683,
32'sd975, 32'sd1511, 32'sd490, 32'sd619, 32'sd1824, 32'sd479,
32'sd978, 32'sd538, 32'sd758, 32'sd509, 32'sd939, 32'sd1507,
32'sd191, 32'sd1371, 32'sd1188, 32'sd1791, 32'sd529, 32'sd1687,
32'sd1773, 32'sd468, 32'sd1221, 32'sd396, 32'sd768, 32'sd1293,
32'sd1411, 32'sd1702, 32'sd591, 32'sd385, 32'sd132, 32'sd1505,
32'sd1861, 32'sd1720, 32'sd1504, 32'sd514, 32'sd294, 32'sd1435,
32'sd531, 32'sd193, 32'sd250, 32'sd1593, 32'sd561, 32'sd462,
32'sd431, 32'sd599, 32'sd910, 32'sd1582, 32'sd646, 32'sd176,
32'sd1879, 32'sd1721, 32'sd1020, 32'sd1192, 32'sd1277, 32'sd1571,
32'sd1527, 32'sd582, 32'sd1881, 32'sd766, 32'sd620, 32'sd1981,
32'sd105, 32'sd183, 32'sd1057, 32'sd328, 32'sd1853, 32'sd994,
32'sd1285, 32'sd1488, 32'sd819, 32'sd1665, 32'sd1536, 32'sd772,
32'sd477, 32'sd443, 32'sd758, 32'sd637, 32'sd764, 32'sd608,
32'sd603, 32'sd597, 32'sd473, 32'sd1805, 32'sd912, 32'sd957,
32'sd1519, 32'sd859, 32'sd1606, 32'sd1824, 32'sd1206, 32'sd1898,
32'sd1587, 32'sd725, 32'sd800, 32'sd952, 32'sd518, 32'sd548,
32'sd1229, 32'sd1740, 32'sd1857, 32'sd1875, 32'sd184, 32'sd467,
32'sd1804, 32'sd850, 32'sd1589, 32'sd1550, 32'sd1983, 32'sd443,
32'sd1704, 32'sd1778, 32'sd1528, 32'sd294, 32'sd440, 32'sd241,
32'sd830, 32'sd395, 32'sd224, 32'sd274, 32'sd1403, 32'sd1396,
32'sd1980, 32'sd1210, 32'sd1617, 32'sd114, 32'sd1943, 32'sd241,
32'sd1877, 32'sd598, 32'sd997, 32'sd676, 32'sd1634, 32'sd377,
32'sd1113, 32'sd1686, 32'sd1794, 32'sd250, 32'sd858, 32'sd1861,
32'sd1516, 32'sd387, 32'sd614, 32'sd1173, 32'sd303, 32'sd1549,
32'sd1099, 32'sd1534, 32'sd657, 32'sd643, 32'sd456, 32'sd659,
32'sd1684, 32'sd619, 32'sd1299, 32'sd352, 32'sd1776, 32'sd1531,
32'sd1184, 32'sd145, 32'sd283, 32'sd778, 32'sd201, 32'sd1321,
32'sd212, 32'sd345, 32'sd1345, 32'sd1589, 32'sd1339, 32'sd392,
32'sd1381, 32'sd440, 32'sd498, 32'sd1187, 32'sd636, 32'sd1579,
32'sd1323, 32'sd1343, 32'sd537, 32'sd862, 32'sd1867, 32'sd797,
32'sd1875, 32'sd865, 32'sd1578, 32'sd446, 32'sd836, 32'sd1460,
32'sd365, 32'sd943, 32'sd753, 32'sd597, 32'sd867, 32'sd1393,
32'sd1792, 32'sd703, 32'sd956, 32'sd1703, 32'sd446, 32'sd593,
32'sd1533, 32'sd116, 32'sd1469, 32'sd821, 32'sd835, 32'sd1056,
32'sd718, 32'sd719, 32'sd1561, 32'sd1009, 32'sd1773, 32'sd523,
32'sd1831, 32'sd846, 32'sd947, 32'sd1590, 32'sd1041, 32'sd1263,
32'sd135, 32'sd1936, 32'sd1589, 32'sd587, 32'sd906, 32'sd345,
32'sd516, 32'sd1314, 32'sd1764, 32'sd703, 32'sd228, 32'sd266,
32'sd1588, 32'sd911, 32'sd1245, 32'sd575, 32'sd1112, 32'sd760,
32'sd1906, 32'sd1733, 32'sd1495, 32'sd802, 32'sd1416, 32'sd1442,
32'sd1177, 32'sd417, 32'sd160, 32'sd420, 32'sd1141, 32'sd1478,
32'sd1136, 32'sd380, 32'sd592, 32'sd1199, 32'sd208, 32'sd1837,
32'sd1793, 32'sd116, 32'sd858, 32'sd388, 32'sd1586, 32'sd465,
32'sd801, 32'sd1666, 32'sd1296, 32'sd755, 32'sd1655, 32'sd1816,
32'sd1292, 32'sd878, 32'sd1262, 32'sd1656, 32'sd1770, 32'sd848,
32'sd781, 32'sd874, 32'sd439, 32'sd878, 32'sd1479, 32'sd1707,
32'sd615, 32'sd581, 32'sd285, 32'sd110, 32'sd126, 32'sd1612,
32'sd374, 32'sd261, 32'sd1865, 32'sd1072, 32'sd1960, 32'sd398,
32'sd1887, 32'sd1462, 32'sd1126, 32'sd745, 32'sd524, 32'sd1084,
32'sd308, 32'sd1077, 32'sd1420, 32'sd542, 32'sd155, 32'sd1797,
32'sd921, 32'sd551, 32'sd1335, 32'sd881, 32'sd377, 32'sd779,
32'sd1697, 32'sd765, 32'sd849, 32'sd382, 32'sd310, 32'sd1449,
32'sd485, 32'sd824, 32'sd1084, 32'sd719, 32'sd1400, 32'sd383,
32'sd724, 32'sd1227, 32'sd1010, 32'sd1866, 32'sd640, 32'sd340,
32'sd1127, 32'sd1723, 32'sd960, 32'sd1153, 32'sd169, 32'sd343,
32'sd1205, 32'sd275, 32'sd1453, 32'sd1343, 32'sd1870, 32'sd652,
32'sd801, 32'sd1932, 32'sd1002, 32'sd899, 32'sd1235, 32'sd1300,
32'sd526, 32'sd440, 32'sd1774, 32'sd934, 32'sd1984, 32'sd1919,
32'sd238, 32'sd496, 32'sd269, 32'sd202, 32'sd1149, 32'sd1863,
32'sd1673, 32'sd1787, 32'sd1070, 32'sd1629, 32'sd281, 32'sd787,
32'sd1626, 32'sd1624, 32'sd609, 32'sd869, 32'sd1009, 32'sd496,
32'sd762, 32'sd1647, 32'sd816, 32'sd1793, 32'sd1662, 32'sd1138,
32'sd1675, 32'sd853, 32'sd428, 32'sd582, 32'sd234, 32'sd1335,
32'sd1943, 32'sd1616, 32'sd1692, 32'sd381, 32'sd355, 32'sd800,
32'sd1452, 32'sd1472, 32'sd178, 32'sd1452, 32'sd1609, 32'sd1491,
32'sd213, 32'sd1713, 32'sd212, 32'sd415, 32'sd1841, 32'sd959,
32'sd530, 32'sd345, 32'sd767, 32'sd927, 32'sd1706, 32'sd499,
32'sd521, 32'sd1089, 32'sd1972, 32'sd1672, 32'sd741, 32'sd969,
32'sd1361, 32'sd121, 32'sd935, 32'sd770, 32'sd1753, 32'sd1439,
32'sd1509, 32'sd129, 32'sd833, 32'sd611, 32'sd430, 32'sd1413,
32'sd1204, 32'sd1930, 32'sd1025, 32'sd1003, 32'sd115, 32'sd1325,
32'sd1409, 32'sd1463, 32'sd120, 32'sd1827, 32'sd1678, 32'sd1377,
32'sd1934, 32'sd1064, 32'sd1134, 32'sd957, 32'sd1940, 32'sd1199,
32'sd1341, 32'sd1514, 32'sd686, 32'sd934, 32'sd1518, 32'sd1158,
32'sd1180, 32'sd959, 32'sd154, 32'sd100, 32'sd1166, 32'sd587,
32'sd932, 32'sd1365, 32'sd709, 32'sd1594, 32'sd881, 32'sd513,
32'sd1147, 32'sd1020, 32'sd1206, 32'sd1810, 32'sd874, 32'sd781,
32'sd1086, 32'sd1817, 32'sd1312, 32'sd1121, 32'sd1960, 32'sd1221,
32'sd152, 32'sd1360, 32'sd1324, 32'sd450, 32'sd1092, 32'sd1554,
32'sd220, 32'sd565, 32'sd276, 32'sd1506, 32'sd1697, 32'sd1410,
32'sd971, 32'sd1213, 32'sd1846, 32'sd1271, 32'sd1815, 32'sd797,
32'sd1500, 32'sd806, 32'sd1000, 32'sd1094, 32'sd698, 32'sd290,
32'sd1589, 32'sd809, 32'sd1413, 32'sd1120, 32'sd1317, 32'sd513,
32'sd1734, 32'sd606, 32'sd1334, 32'sd1114, 32'sd1275, 32'sd1029,
32'sd1884, 32'sd1521, 32'sd1575, 32'sd1141, 32'sd1533, 32'sd743,
32'sd491, 32'sd1091, 32'sd1621, 32'sd325, 32'sd273, 32'sd373,
32'sd1971, 32'sd666, 32'sd1401, 32'sd1043, 32'sd1685, 32'sd539,
32'sd309, 32'sd600, 32'sd1411, 32'sd508, 32'sd372, 32'sd614,
32'sd1634, 32'sd1372, 32'sd644, 32'sd1810, 32'sd1461, 32'sd612,
32'sd982, 32'sd1312, 32'sd1383, 32'sd1205, 32'sd182, 32'sd1652,
32'sd645, 32'sd971, 32'sd596, 32'sd546, 32'sd314, 32'sd1784,
32'sd1337, 32'sd1943, 32'sd782, 32'sd1313, 32'sd362, 32'sd991,
32'sd1280, 32'sd1028, 32'sd143, 32'sd552, 32'sd615, 32'sd1120,
32'sd400, 32'sd1225, 32'sd482, 32'sd1756, 32'sd1430, 32'sd1186,
32'sd731, 32'sd1582, 32'sd648, 32'sd1051, 32'sd556, 32'sd211,
32'sd1603, 32'sd1775, 32'sd1484, 32'sd1536, 32'sd1732, 32'sd577,
32'sd1714, 32'sd746, 32'sd1464, 32'sd1183, 32'sd1415, 32'sd1165,
32'sd1248, 32'sd1467, 32'sd1440, 32'sd526, 32'sd509, 32'sd1755,
32'sd1234, 32'sd1965, 32'sd1058, 32'sd1688, 32'sd1886, 32'sd915,
32'sd1532, 32'sd457, 32'sd138, 32'sd1786, 32'sd597, 32'sd1279,
32'sd351, 32'sd412, 32'sd1124, 32'sd1975, 32'sd1407, 32'sd837,
32'sd168, 32'sd338, 32'sd599, 32'sd1623, 32'sd684, 32'sd330,
32'sd300, 32'sd1336, 32'sd1438, 32'sd1211, 32'sd874, 32'sd727,
32'sd1465, 32'sd1269, 32'sd1458, 32'sd1468, 32'sd596, 32'sd1559,
32'sd1454, 32'sd1465, 32'sd1380, 32'sd1658, 32'sd1453, 32'sd1438,
32'sd1275, 32'sd975, 32'sd329, 32'sd637, 32'sd1054, 32'sd1146,
32'sd1124, 32'sd188, 32'sd211, 32'sd1472, 32'sd298, 32'sd1192,
32'sd960, 32'sd1228, 32'sd478, 32'sd1666, 32'sd214, 32'sd445,
32'sd888, 32'sd360, 32'sd873, 32'sd1749, 32'sd1581, 32'sd824,
32'sd1453, 32'sd403, 32'sd679, 32'sd1681, 32'sd1884, 32'sd1560,
32'sd1406, 32'sd1006, 32'sd874, 32'sd183, 32'sd334, 32'sd849,
32'sd1731, 32'sd963, 32'sd881, 32'sd1060, 32'sd1240, 32'sd1775,
32'sd480, 32'sd1204, 32'sd1977, 32'sd1252, 32'sd575, 32'sd303,
32'sd123, 32'sd1951, 32'sd1945, 32'sd1166, 32'sd473, 32'sd401,
32'sd931, 32'sd981, 32'sd1765, 32'sd1771, 32'sd1674, 32'sd1656,
32'sd1739, 32'sd198, 32'sd1339, 32'sd704, 32'sd316, 32'sd1999,
32'sd641, 32'sd402, 32'sd994, 32'sd1198, 32'sd1964, 32'sd1240,
32'sd283, 32'sd1982, 32'sd381, 32'sd404, 32'sd1797, 32'sd1602,
32'sd1888, 32'sd305, 32'sd1581, 32'sd1798, 32'sd1312, 32'sd1784,
32'sd1818, 32'sd152, 32'sd895, 32'sd102, 32'sd863, 32'sd497,
32'sd1567, 32'sd195, 32'sd746, 32'sd1016, 32'sd862, 32'sd1704,
32'sd1696, 32'sd418, 32'sd858, 32'sd538, 32'sd1583, 32'sd1507,
32'sd1065, 32'sd1028, 32'sd777, 32'sd238, 32'sd458, 32'sd1319,
32'sd466, 32'sd1332, 32'sd164, 32'sd1538, 32'sd837, 32'sd1484,
32'sd1052, 32'sd1093, 32'sd1267, 32'sd1143, 32'sd1699, 32'sd1110,
32'sd1143, 32'sd1869, 32'sd1187, 32'sd455, 32'sd898, 32'sd1664,
32'sd1508, 32'sd1240, 32'sd1591, 32'sd1446, 32'sd422, 32'sd1636,
32'sd1781, 32'sd622, 32'sd579, 32'sd1165, 32'sd1809, 32'sd1510,
32'sd1614, 32'sd1871, 32'sd674, 32'sd1249, 32'sd422, 32'sd847,
32'sd1731, 32'sd341, 32'sd1868, 32'sd1928, 32'sd333, 32'sd337,
32'sd1496, 32'sd638, 32'sd437, 32'sd916, 32'sd594, 32'sd303,
32'sd1273, 32'sd660, 32'sd1584, 32'sd852, 32'sd978, 32'sd1337,
32'sd1637, 32'sd338, 32'sd743, 32'sd1389, 32'sd402, 32'sd1462,
32'sd1252, 32'sd1614, 32'sd1375, 32'sd1411, 32'sd387, 32'sd862,
32'sd593, 32'sd1744, 32'sd494, 32'sd540, 32'sd643, 32'sd1280,
32'sd1613, 32'sd587, 32'sd1698, 32'sd712, 32'sd1335, 32'sd1986,
32'sd1618, 32'sd1720, 32'sd1222, 32'sd794, 32'sd896, 32'sd1674,
32'sd1186, 32'sd1092, 32'sd591, 32'sd519, 32'sd137, 32'sd319,
32'sd994, 32'sd695, 32'sd952, 32'sd710, 32'sd1572, 32'sd812,
32'sd1583, 32'sd1793, 32'sd673, 32'sd1777, 32'sd954, 32'sd1504,
32'sd1536, 32'sd279, 32'sd895, 32'sd1296, 32'sd148, 32'sd462,
32'sd1341, 32'sd1970, 32'sd1950, 32'sd1588, 32'sd258, 32'sd673,
32'sd1775, 32'sd1838, 32'sd281, 32'sd677, 32'sd703, 32'sd708,
32'sd205, 32'sd1259, 32'sd893, 32'sd1025, 32'sd411, 32'sd941,
32'sd1855, 32'sd744, 32'sd1666, 32'sd1372, 32'sd1660, 32'sd1877,
32'sd713, 32'sd132, 32'sd432, 32'sd378, 32'sd118, 32'sd1547,
32'sd1182, 32'sd1143, 32'sd358, 32'sd1138, 32'sd742, 32'sd798,
32'sd1034, 32'sd279, 32'sd515, 32'sd465, 32'sd447, 32'sd552,
32'sd1779, 32'sd1848, 32'sd1924, 32'sd1346, 32'sd1427, 32'sd497,
32'sd644, 32'sd1630, 32'sd1087, 32'sd1483, 32'sd1609, 32'sd263,
32'sd880, 32'sd1676, 32'sd505, 32'sd890, 32'sd1239, 32'sd626,
32'sd921, 32'sd1654, 32'sd301, 32'sd1507, 32'sd1578, 32'sd1352,
32'sd1678, 32'sd622, 32'sd1874, 32'sd1886, 32'sd383, 32'sd1705,
32'sd698, 32'sd1273, 32'sd340, 32'sd600, 32'sd1314, 32'sd1574,
32'sd921, 32'sd297, 32'sd1615, 32'sd642, 32'sd515, 32'sd568,
32'sd647, 32'sd1650, 32'sd1524, 32'sd1340, 32'sd1320, 32'sd1207,
32'sd143, 32'sd512, 32'sd469, 32'sd785, 32'sd1827, 32'sd1308,
32'sd1785, 32'sd200, 32'sd155, 32'sd886, 32'sd1578, 32'sd1041,
32'sd523, 32'sd1438, 32'sd1795, 32'sd542, 32'sd933, 32'sd1281,
32'sd1613, 32'sd1917, 32'sd1215, 32'sd924, 32'sd986, 32'sd1806,
32'sd1926, 32'sd1546, 32'sd1549, 32'sd931, 32'sd1083, 32'sd1786,
32'sd1993, 32'sd447, 32'sd976, 32'sd1856, 32'sd1937, 32'sd1080,
32'sd1301, 32'sd1735, 32'sd274, 32'sd1309, 32'sd234, 32'sd1979,
32'sd307, 32'sd949, 32'sd1219, 32'sd571, 32'sd1721, 32'sd542,
32'sd849, 32'sd1768, 32'sd574, 32'sd1817, 32'sd543, 32'sd125,
32'sd899, 32'sd1695, 32'sd1263, 32'sd423, 32'sd850, 32'sd467,
32'sd240, 32'sd140, 32'sd1554, 32'sd1987, 32'sd1666, 32'sd1796,
32'sd1114, 32'sd985, 32'sd374, 32'sd1735, 32'sd1034, 32'sd567,
32'sd524, 32'sd769, 32'sd208, 32'sd566, 32'sd1375, 32'sd1955,
32'sd434, 32'sd882, 32'sd217, 32'sd377, 32'sd1716, 32'sd1154,
32'sd1248, 32'sd1060, 32'sd878, 32'sd1874, 32'sd1934, 32'sd1602,
32'sd1051, 32'sd431, 32'sd404, 32'sd1492, 32'sd1308, 32'sd120,
32'sd1317, 32'sd559, 32'sd805, 32'sd829, 32'sd868, 32'sd887,
32'sd496, 32'sd972, 32'sd423, 32'sd1835, 32'sd1389, 32'sd1295,
32'sd1758, 32'sd1201, 32'sd885, 32'sd1217, 32'sd1352, 32'sd1686,
32'sd1249, 32'sd1903, 32'sd845, 32'sd1925, 32'sd1682, 32'sd1273,
32'sd1255, 32'sd1041, 32'sd180, 32'sd1992, 32'sd1701, 32'sd937,
32'sd1638, 32'sd880, 32'sd1736, 32'sd366, 32'sd656, 32'sd274,
32'sd1133, 32'sd1789, 32'sd503, 32'sd1650, 32'sd1681, 32'sd530,
32'sd1953, 32'sd196, 32'sd1273, 32'sd1652, 32'sd1222, 32'sd1339,
32'sd1414, 32'sd644, 32'sd1582, 32'sd1001, 32'sd1818, 32'sd583,
32'sd1071, 32'sd1028, 32'sd652, 32'sd422, 32'sd455, 32'sd1678,
32'sd427, 32'sd401, 32'sd806, 32'sd1486, 32'sd686, 32'sd604,
32'sd1638, 32'sd470, 32'sd378, 32'sd1538, 32'sd1029, 32'sd337,
32'sd391, 32'sd1471, 32'sd491, 32'sd425, 32'sd121, 32'sd1299,
32'sd1133, 32'sd195, 32'sd1770, 32'sd365, 32'sd820, 32'sd674,
32'sd1276, 32'sd1579, 32'sd879, 32'sd1538, 32'sd1131, 32'sd227,
32'sd201, 32'sd1167, 32'sd743, 32'sd486, 32'sd746, 32'sd1185,
32'sd1007, 32'sd613, 32'sd1192, 32'sd1924, 32'sd1582, 32'sd411,
32'sd1531, 32'sd187, 32'sd139, 32'sd1306, 32'sd122, 32'sd238,
32'sd109, 32'sd871, 32'sd1273, 32'sd180, 32'sd471, 32'sd1355,
32'sd147, 32'sd767, 32'sd707, 32'sd200, 32'sd435, 32'sd422,
32'sd856, 32'sd1548, 32'sd1845, 32'sd1555, 32'sd1038, 32'sd730,
32'sd1275, 32'sd1861, 32'sd1398, 32'sd318, 32'sd1307, 32'sd1505,
32'sd1461, 32'sd106, 32'sd1562, 32'sd717, 32'sd695, 32'sd1049,
32'sd1228, 32'sd1705, 32'sd1940, 32'sd1172, 32'sd1968, 32'sd1488,
32'sd1249, 32'sd1735, 32'sd1070, 32'sd1858, 32'sd566, 32'sd488,
32'sd1608, 32'sd474, 32'sd402, 32'sd885, 32'sd1467, 32'sd1548,
32'sd1799, 32'sd982, 32'sd266, 32'sd1466, 32'sd105, 32'sd1925,
32'sd1297, 32'sd871, 32'sd182, 32'sd1713, 32'sd1371, 32'sd283,
32'sd1456, 32'sd1323, 32'sd633, 32'sd1908, 32'sd1453, 32'sd1636,
32'sd1221, 32'sd1362, 32'sd1720, 32'sd1730, 32'sd1327, 32'sd1231,
32'sd758, 32'sd1886, 32'sd1011, 32'sd1070, 32'sd1465, 32'sd1903,
32'sd1813, 32'sd431, 32'sd1413, 32'sd895, 32'sd1844, 32'sd184,
32'sd421, 32'sd1099, 32'sd1230, 32'sd1027, 32'sd1976, 32'sd122,
32'sd107, 32'sd974, 32'sd313, 32'sd482, 32'sd154, 32'sd503,
32'sd737, 32'sd775, 32'sd593, 32'sd1384, 32'sd298, 32'sd412,
32'sd432, 32'sd1343, 32'sd505, 32'sd105, 32'sd1274, 32'sd980,
32'sd1351, 32'sd384, 32'sd1297, 32'sd192, 32'sd954, 32'sd855,
32'sd1610, 32'sd759, 32'sd288, 32'sd1276, 32'sd860, 32'sd1349,
32'sd1891, 32'sd1774, 32'sd1853, 32'sd350, 32'sd1661, 32'sd1095,
32'sd1370, 32'sd1575, 32'sd340, 32'sd1535, 32'sd980, 32'sd1357,
32'sd360, 32'sd892, 32'sd350, 32'sd494, 32'sd727, 32'sd235,
32'sd1050, 32'sd793, 32'sd1177, 32'sd1859, 32'sd1234, 32'sd133,
32'sd578, 32'sd282, 32'sd1493, 32'sd180, 32'sd1909, 32'sd1165,
32'sd1568, 32'sd869, 32'sd1908, 32'sd742, 32'sd556, 32'sd1403,
32'sd1109, 32'sd1176, 32'sd920, 32'sd1894, 32'sd1437, 32'sd1745,
32'sd1037, 32'sd891, 32'sd1712, 32'sd952, 32'sd947, 32'sd958,
32'sd207, 32'sd1066, 32'sd565, 32'sd1108, 32'sd1620, 32'sd1999,
32'sd1385, 32'sd1028, 32'sd776, 32'sd1130, 32'sd1845, 32'sd972,
32'sd1662, 32'sd427, 32'sd1345, 32'sd112, 32'sd1815, 32'sd563,
32'sd1204, 32'sd643, 32'sd1742, 32'sd1108, 32'sd764, 32'sd1978,
32'sd533, 32'sd458, 32'sd354, 32'sd1624, 32'sd304, 32'sd1918,
32'sd433, 32'sd122, 32'sd1643, 32'sd700, 32'sd228, 32'sd1560,
32'sd873, 32'sd1954, 32'sd260, 32'sd733, 32'sd1891, 32'sd1798,
32'sd661, 32'sd442, 32'sd1781, 32'sd1807, 32'sd1311, 32'sd1099,
32'sd105, 32'sd1349, 32'sd1546, 32'sd396, 32'sd1408, 32'sd1360,
32'sd1016, 32'sd1037, 32'sd1814, 32'sd320, 32'sd1510, 32'sd1314,
32'sd1115, 32'sd1335, 32'sd830, 32'sd1062, 32'sd825, 32'sd1864,
32'sd472, 32'sd1643, 32'sd744, 32'sd724, 32'sd772, 32'sd1025,
32'sd1235, 32'sd633, 32'sd585, 32'sd346, 32'sd1572, 32'sd1244,
32'sd1687, 32'sd1807, 32'sd940, 32'sd1565, 32'sd1062, 32'sd112,
32'sd810, 32'sd1407, 32'sd1195, 32'sd445, 32'sd1316, 32'sd1563,
32'sd1200, 32'sd1032, 32'sd388, 32'sd1748, 32'sd1070, 32'sd911,
32'sd633, 32'sd354, 32'sd945, 32'sd1376, 32'sd838, 32'sd1996,
32'sd1735, 32'sd1492, 32'sd1098, 32'sd932, 32'sd803, 32'sd1372,
32'sd1871, 32'sd634, 32'sd1660, 32'sd1678, 32'sd1718, 32'sd784,
32'sd1319, 32'sd1266, 32'sd961, 32'sd240, 32'sd501, 32'sd1949,
32'sd1871, 32'sd898, 32'sd985, 32'sd504, 32'sd289, 32'sd1532,
32'sd828, 32'sd1134, 32'sd1044, 32'sd1053, 32'sd757, 32'sd795,
32'sd1684, 32'sd940, 32'sd1338, 32'sd163, 32'sd1755, 32'sd1072,
32'sd1406, 32'sd1995, 32'sd177, 32'sd1036, 32'sd556, 32'sd400,
32'sd847, 32'sd1228, 32'sd654, 32'sd1647, 32'sd1876, 32'sd1961,
32'sd779, 32'sd1866, 32'sd818, 32'sd1162, 32'sd1211, 32'sd1914,
32'sd1693, 32'sd1365, 32'sd494, 32'sd292, 32'sd1978, 32'sd1818,
32'sd927, 32'sd1303, 32'sd1460, 32'sd1050, 32'sd1890, 32'sd1175,
32'sd1286, 32'sd439, 32'sd1179, 32'sd205, 32'sd977, 32'sd168,
32'sd1425, 32'sd600, 32'sd1214, 32'sd736, 32'sd1155, 32'sd1333,
32'sd1730, 32'sd866, 32'sd1404, 32'sd384, 32'sd1277, 32'sd1042,
32'sd1105, 32'sd879, 32'sd194, 32'sd136, 32'sd1038, 32'sd1476,
32'sd1480, 32'sd1143, 32'sd260, 32'sd1667, 32'sd214, 32'sd1534,
32'sd668, 32'sd122, 32'sd1062, 32'sd1029, 32'sd1629, 32'sd770,
32'sd1175, 32'sd927, 32'sd1796, 32'sd1572, 32'sd1454, 32'sd1449,
32'sd1500, 32'sd1008, 32'sd497, 32'sd496, 32'sd1960, 32'sd436,
32'sd1783, 32'sd464, 32'sd982, 32'sd1606, 32'sd644, 32'sd270,
32'sd583, 32'sd705, 32'sd1680, 32'sd1532, 32'sd244, 32'sd161,
32'sd1366, 32'sd1172, 32'sd1295, 32'sd1200, 32'sd529, 32'sd991,
32'sd225, 32'sd1791, 32'sd121, 32'sd1316, 32'sd1439, 32'sd304,
32'sd1757, 32'sd1726, 32'sd1231, 32'sd747, 32'sd344, 32'sd1446,
32'sd132, 32'sd1104, 32'sd473, 32'sd1291, 32'sd469, 32'sd605,
32'sd487, 32'sd1214, 32'sd1137, 32'sd1846, 32'sd1514, 32'sd114,
32'sd601, 32'sd1817, 32'sd513, 32'sd1160, 32'sd1453, 32'sd1603,
32'sd892, 32'sd869, 32'sd1036, 32'sd495, 32'sd751, 32'sd412,
32'sd157, 32'sd1986, 32'sd195, 32'sd383, 32'sd1321, 32'sd153,
32'sd724, 32'sd211, 32'sd647, 32'sd617, 32'sd627, 32'sd1813,
32'sd1358, 32'sd1757, 32'sd1690, 32'sd1692, 32'sd1523, 32'sd312,
32'sd441, 32'sd642, 32'sd1169, 32'sd735, 32'sd945, 32'sd389,
32'sd566, 32'sd968, 32'sd1711, 32'sd105, 32'sd740, 32'sd1560,
32'sd1489, 32'sd269, 32'sd115, 32'sd1240, 32'sd413, 32'sd275,
32'sd666, 32'sd684, 32'sd471, 32'sd1440, 32'sd1666, 32'sd135,
32'sd884, 32'sd944, 32'sd1502, 32'sd449, 32'sd781, 32'sd1817,
32'sd664, 32'sd135, 32'sd1842, 32'sd439, 32'sd669, 32'sd1889,
32'sd1875, 32'sd1742, 32'sd239, 32'sd267, 32'sd1086, 32'sd1807,
32'sd1261, 32'sd673, 32'sd1695, 32'sd1422, 32'sd1104, 32'sd319,
32'sd610, 32'sd1610, 32'sd285, 32'sd614, 32'sd989, 32'sd1723,
32'sd1617, 32'sd199, 32'sd628, 32'sd438, 32'sd236, 32'sd806,
32'sd1275, 32'sd199, 32'sd1975, 32'sd1149, 32'sd1798, 32'sd1241,
32'sd1169, 32'sd1323, 32'sd1248, 32'sd1994, 32'sd152, 32'sd855,
32'sd1397, 32'sd523, 32'sd1740, 32'sd1625, 32'sd1381, 32'sd537,
32'sd1519, 32'sd869, 32'sd1500, 32'sd1650, 32'sd212, 32'sd803,
32'sd375, 32'sd919, 32'sd1827, 32'sd1925, 32'sd703, 32'sd636,
32'sd1504, 32'sd1188, 32'sd897, 32'sd1642, 32'sd1073, 32'sd164,
32'sd455, 32'sd1088, 32'sd574, 32'sd1455, 32'sd732, 32'sd1409,
32'sd1999, 32'sd1949, 32'sd1679, 32'sd1940, 32'sd141, 32'sd1519,
32'sd820, 32'sd179, 32'sd402, 32'sd1892, 32'sd1402, 32'sd796,
32'sd971, 32'sd370, 32'sd751, 32'sd1095, 32'sd1558, 32'sd672,
32'sd248, 32'sd1608, 32'sd858, 32'sd1189, 32'sd1482, 32'sd759,
32'sd719, 32'sd237, 32'sd628, 32'sd1858, 32'sd668, 32'sd1057,
32'sd1478, 32'sd854, 32'sd379, 32'sd1026, 32'sd1071, 32'sd201,
32'sd1930, 32'sd548, 32'sd1955, 32'sd242, 32'sd305, 32'sd692,
32'sd155, 32'sd1996, 32'sd1542, 32'sd984, 32'sd209, 32'sd373,
32'sd1504, 32'sd1101, 32'sd1337, 32'sd494, 32'sd1337, 32'sd110,
32'sd1178, 32'sd1173, 32'sd753, 32'sd751, 32'sd845, 32'sd1984,
32'sd442, 32'sd587, 32'sd853, 32'sd1553, 32'sd726, 32'sd1330,
32'sd142, 32'sd1287, 32'sd1729, 32'sd1891, 32'sd127, 32'sd1251,
32'sd1706, 32'sd1045, 32'sd847, 32'sd1799, 32'sd567, 32'sd795,
32'sd1975, 32'sd570, 32'sd986, 32'sd1049, 32'sd1833, 32'sd973,
32'sd1337, 32'sd1810, 32'sd521, 32'sd215, 32'sd336, 32'sd1261,
32'sd1420, 32'sd1387, 32'sd287, 32'sd433, 32'sd1035, 32'sd585,
32'sd498, 32'sd1384, 32'sd615, 32'sd1158, 32'sd1443, 32'sd1144,
32'sd1736, 32'sd837, 32'sd108, 32'sd313, 32'sd1870, 32'sd1634,
32'sd1808, 32'sd974, 32'sd1748, 32'sd1412, 32'sd998, 32'sd652,
32'sd704, 32'sd357, 32'sd769, 32'sd1732, 32'sd582, 32'sd792,
32'sd126, 32'sd1546, 32'sd590, 32'sd1563, 32'sd1371, 32'sd502,
32'sd1525, 32'sd1476, 32'sd611, 32'sd678, 32'sd638, 32'sd1789,
32'sd346, 32'sd1980, 32'sd797, 32'sd1837, 32'sd953, 32'sd895,
32'sd1357, 32'sd484, 32'sd619, 32'sd1824, 32'sd1523, 32'sd475,
32'sd983, 32'sd766, 32'sd1724, 32'sd273, 32'sd1900, 32'sd157,
32'sd1233, 32'sd1147, 32'sd1935, 32'sd242, 32'sd1487, 32'sd527,
32'sd625, 32'sd1229, 32'sd1512, 32'sd1915, 32'sd1009, 32'sd482,
32'sd1992, 32'sd1542, 32'sd254, 32'sd824, 32'sd1579, 32'sd963,
32'sd909, 32'sd560, 32'sd1286, 32'sd1989, 32'sd1599, 32'sd818,
32'sd1838, 32'sd371, 32'sd1558, 32'sd1036, 32'sd808, 32'sd1569,
32'sd316, 32'sd597, 32'sd173, 32'sd1713, 32'sd1766, 32'sd1603,
32'sd1812, 32'sd447, 32'sd1642, 32'sd232, 32'sd1102, 32'sd1500,
32'sd249, 32'sd1384, 32'sd1308, 32'sd540, 32'sd1087, 32'sd1207,
32'sd184, 32'sd277, 32'sd683, 32'sd972, 32'sd1767, 32'sd773,
32'sd577, 32'sd1868, 32'sd370, 32'sd1909, 32'sd1801, 32'sd1568,
32'sd1440, 32'sd307, 32'sd1961, 32'sd1015, 32'sd299, 32'sd416,
32'sd696, 32'sd671, 32'sd1868, 32'sd278, 32'sd1970, 32'sd667,
32'sd178, 32'sd1825, 32'sd698, 32'sd434, 32'sd1985, 32'sd1732,
32'sd587, 32'sd938, 32'sd1260, 32'sd832, 32'sd410, 32'sd1572,
32'sd1798, 32'sd847, 32'sd1527, 32'sd242, 32'sd1327, 32'sd1834,
32'sd1450, 32'sd1936, 32'sd1849, 32'sd848, 32'sd468, 32'sd349,
32'sd1483, 32'sd578, 32'sd120, 32'sd466, 32'sd1885, 32'sd243,
32'sd328, 32'sd1391, 32'sd274, 32'sd1362, 32'sd1939, 32'sd1031,
32'sd559, 32'sd781, 32'sd450, 32'sd1158, 32'sd113, 32'sd1396,
32'sd1610, 32'sd1847, 32'sd730, 32'sd366, 32'sd1639, 32'sd1956,
32'sd1477, 32'sd576, 32'sd1434, 32'sd907, 32'sd1465, 32'sd230,
32'sd467, 32'sd277, 32'sd866, 32'sd1149, 32'sd1883, 32'sd1313,
32'sd1231, 32'sd1571, 32'sd409, 32'sd348, 32'sd699, 32'sd571,
32'sd932, 32'sd539, 32'sd633, 32'sd1574, 32'sd838, 32'sd1622,
32'sd267, 32'sd329, 32'sd1181, 32'sd1717, 32'sd1353, 32'sd1680,
32'sd1569, 32'sd509, 32'sd281, 32'sd848, 32'sd619, 32'sd1308,
32'sd349, 32'sd487, 32'sd1445, 32'sd1307, 32'sd1102, 32'sd218,
32'sd1931, 32'sd249, 32'sd1375, 32'sd556, 32'sd1008, 32'sd1494,
32'sd405, 32'sd1001, 32'sd933, 32'sd994, 32'sd1763, 32'sd1095,
32'sd569, 32'sd1469, 32'sd999, 32'sd491, 32'sd1135, 32'sd1009,
32'sd849, 32'sd126, 32'sd947, 32'sd1731, 32'sd1974, 32'sd774,
32'sd659, 32'sd1958, 32'sd1039, 32'sd1460, 32'sd1934, 32'sd1027,
32'sd1061, 32'sd244, 32'sd153, 32'sd1364, 32'sd661, 32'sd1857,
32'sd968, 32'sd419, 32'sd1493, 32'sd1765, 32'sd1967, 32'sd1434,
32'sd1444, 32'sd1523, 32'sd1692, 32'sd422, 32'sd131, 32'sd720,
32'sd429, 32'sd320, 32'sd633, 32'sd1374, 32'sd1034, 32'sd1491,
32'sd132, 32'sd165, 32'sd1087, 32'sd282, 32'sd1257, 32'sd206,
32'sd173, 32'sd539, 32'sd1517, 32'sd842, 32'sd1711, 32'sd1684,
32'sd1329, 32'sd1557, 32'sd808, 32'sd1596, 32'sd139, 32'sd690,
32'sd1566, 32'sd699, 32'sd961, 32'sd261, 32'sd1762, 32'sd1350,
32'sd356, 32'sd1927, 32'sd756, 32'sd1850, 32'sd1002, 32'sd251,
32'sd578, 32'sd1119, 32'sd276, 32'sd1031, 32'sd1365, 32'sd564,
32'sd147, 32'sd1474, 32'sd472, 32'sd680, 32'sd1483, 32'sd321,
32'sd321, 32'sd635, 32'sd501, 32'sd1473, 32'sd1361, 32'sd563,
32'sd1970, 32'sd1425, 32'sd1415, 32'sd506, 32'sd610, 32'sd231,
32'sd1899, 32'sd1927, 32'sd443, 32'sd842, 32'sd562, 32'sd1384,
32'sd620, 32'sd1994, 32'sd476, 32'sd845, 32'sd508, 32'sd854,
32'sd1153, 32'sd1500, 32'sd519, 32'sd1412, 32'sd969, 32'sd1227,
32'sd1401, 32'sd1499, 32'sd1505, 32'sd1789, 32'sd393, 32'sd339,
32'sd224, 32'sd1438, 32'sd826, 32'sd1813, 32'sd370, 32'sd181,
32'sd594, 32'sd856, 32'sd1662, 32'sd906, 32'sd810, 32'sd476,
32'sd231, 32'sd762, 32'sd1409, 32'sd1417, 32'sd1328, 32'sd1541,
32'sd1110, 32'sd968, 32'sd1179, 32'sd688, 32'sd1251, 32'sd741,
32'sd1144, 32'sd1098, 32'sd238, 32'sd1323, 32'sd361, 32'sd863,
32'sd792, 32'sd1767, 32'sd686, 32'sd1230, 32'sd1899, 32'sd1777,
32'sd1023, 32'sd1565, 32'sd904, 32'sd1206, 32'sd554, 32'sd776,
32'sd178, 32'sd1502, 32'sd825, 32'sd1987, 32'sd622, 32'sd1032,
32'sd464, 32'sd663, 32'sd581, 32'sd168, 32'sd1928, 32'sd908,
32'sd1806, 32'sd282, 32'sd1396, 32'sd1136, 32'sd732, 32'sd967,
32'sd292, 32'sd184, 32'sd1652, 32'sd134, 32'sd613, 32'sd1723,
32'sd1655, 32'sd594, 32'sd930, 32'sd1881, 32'sd354, 32'sd1017,
32'sd1291, 32'sd950, 32'sd1044, 32'sd688, 32'sd1971, 32'sd759,
32'sd1853, 32'sd1405, 32'sd897, 32'sd235, 32'sd430, 32'sd847,
32'sd1614, 32'sd233, 32'sd625, 32'sd1050, 32'sd1655, 32'sd1143,
32'sd1595, 32'sd1823, 32'sd1546, 32'sd720, 32'sd608, 32'sd643,
32'sd1943, 32'sd1286, 32'sd169, 32'sd1084, 32'sd1481, 32'sd1108,
32'sd635, 32'sd315, 32'sd1841, 32'sd621, 32'sd1376, 32'sd1720,
32'sd1901, 32'sd1606, 32'sd660, 32'sd1820, 32'sd916, 32'sd1926,
32'sd1162, 32'sd1452, 32'sd345, 32'sd984, 32'sd585, 32'sd1049,
32'sd1027, 32'sd1611, 32'sd855, 32'sd1273, 32'sd1719, 32'sd1629,
32'sd1827, 32'sd143, 32'sd1197, 32'sd833, 32'sd854, 32'sd1792,
32'sd1860, 32'sd1267, 32'sd1423, 32'sd659, 32'sd1270, 32'sd1843,
32'sd924, 32'sd209, 32'sd1150, 32'sd1656, 32'sd711, 32'sd1715,
32'sd1801, 32'sd1533, 32'sd1514, 32'sd343, 32'sd171, 32'sd1145,
32'sd1373, 32'sd1399, 32'sd479, 32'sd931, 32'sd148, 32'sd935,
32'sd1893, 32'sd1271, 32'sd1818, 32'sd506, 32'sd1228, 32'sd1607,
32'sd1017, 32'sd1477, 32'sd106, 32'sd1566, 32'sd234, 32'sd331,
32'sd781, 32'sd308, 32'sd535, 32'sd1610, 32'sd852, 32'sd1795,
32'sd1831, 32'sd1289, 32'sd154, 32'sd360, 32'sd211, 32'sd218,
32'sd404, 32'sd1371, 32'sd1387, 32'sd1474, 32'sd940, 32'sd160,
32'sd425, 32'sd1992, 32'sd1893, 32'sd1286, 32'sd496, 32'sd165,
32'sd625, 32'sd789, 32'sd1497, 32'sd273, 32'sd315, 32'sd485,
32'sd1055, 32'sd1747, 32'sd430, 32'sd1140, 32'sd1086, 32'sd792,
32'sd1055, 32'sd553, 32'sd224, 32'sd1801, 32'sd1573, 32'sd1508,
32'sd1114, 32'sd829, 32'sd1015, 32'sd880, 32'sd1077, 32'sd662,
32'sd892, 32'sd1756, 32'sd117, 32'sd1981, 32'sd811, 32'sd1865,
32'sd651, 32'sd1776, 32'sd917, 32'sd624, 32'sd170, 32'sd966,
32'sd1037, 32'sd1254, 32'sd1303, 32'sd1773, 32'sd1906, 32'sd818,
32'sd905, 32'sd1762, 32'sd1850, 32'sd821, 32'sd1798, 32'sd914,
32'sd856, 32'sd257, 32'sd514, 32'sd1428, 32'sd1587, 32'sd129,
32'sd1676, 32'sd1477, 32'sd1187, 32'sd593, 32'sd930, 32'sd1676,
32'sd1346, 32'sd143, 32'sd482, 32'sd1564, 32'sd848, 32'sd1775,
32'sd328, 32'sd650, 32'sd1781, 32'sd984, 32'sd1974, 32'sd1425,
32'sd1134, 32'sd1426, 32'sd1759, 32'sd1383, 32'sd776, 32'sd1082,
32'sd1678, 32'sd1046, 32'sd1305, 32'sd1376, 32'sd1814, 32'sd1598,
32'sd902, 32'sd446, 32'sd1662, 32'sd424, 32'sd1048, 32'sd1503,
32'sd1140, 32'sd1127, 32'sd471, 32'sd373, 32'sd566, 32'sd1293,
32'sd1870, 32'sd719, 32'sd1425, 32'sd1644, 32'sd638, 32'sd156,
32'sd1740, 32'sd1362, 32'sd1213, 32'sd849, 32'sd410, 32'sd567,
32'sd561, 32'sd576, 32'sd1009, 32'sd1322, 32'sd459, 32'sd881,
32'sd1074, 32'sd1497, 32'sd680, 32'sd1640, 32'sd300, 32'sd1460,
32'sd1286, 32'sd379, 32'sd762, 32'sd107, 32'sd1726, 32'sd1486,
32'sd1902, 32'sd461, 32'sd1950, 32'sd472, 32'sd835, 32'sd1660,
32'sd611, 32'sd746, 32'sd839, 32'sd1911, 32'sd1776, 32'sd1173,
32'sd1115, 32'sd1059, 32'sd1550, 32'sd971, 32'sd1657, 32'sd1065,
32'sd1562, 32'sd1316, 32'sd739, 32'sd647, 32'sd517, 32'sd1895,
32'sd1377, 32'sd600, 32'sd274, 32'sd592, 32'sd830, 32'sd1706,
32'sd296, 32'sd879, 32'sd1154, 32'sd1792, 32'sd832, 32'sd842,
32'sd1898, 32'sd252, 32'sd1220, 32'sd560, 32'sd1435, 32'sd557,
32'sd711, 32'sd1440, 32'sd1976, 32'sd1655, 32'sd1078, 32'sd404,
32'sd364, 32'sd718, 32'sd1846, 32'sd1996, 32'sd1347, 32'sd1350,
32'sd1393, 32'sd239, 32'sd387, 32'sd695, 32'sd787, 32'sd884,
32'sd798, 32'sd596, 32'sd626, 32'sd1459, 32'sd1771, 32'sd233,
32'sd1900, 32'sd738, 32'sd1313, 32'sd1067, 32'sd335, 32'sd299,
32'sd1364, 32'sd1740, 32'sd435, 32'sd1018, 32'sd1057, 32'sd1858,
32'sd1179, 32'sd1383, 32'sd134, 32'sd932, 32'sd145, 32'sd1795,
32'sd199, 32'sd1679, 32'sd151, 32'sd691, 32'sd242, 32'sd1791,
32'sd1467, 32'sd246, 32'sd503, 32'sd939, 32'sd782, 32'sd291,
32'sd1120, 32'sd1833, 32'sd817, 32'sd687, 32'sd412, 32'sd1300,
32'sd788, 32'sd1750, 32'sd761, 32'sd215, 32'sd1303, 32'sd1719,
32'sd336, 32'sd838, 32'sd1365, 32'sd1775, 32'sd1265, 32'sd1705,
32'sd1256, 32'sd1724, 32'sd1619, 32'sd1528, 32'sd708, 32'sd343,
32'sd718, 32'sd493, 32'sd864, 32'sd312, 32'sd229, 32'sd1781,
32'sd1562, 32'sd598, 32'sd700, 32'sd1125, 32'sd1839, 32'sd1784,
32'sd1753, 32'sd1796, 32'sd1476, 32'sd875, 32'sd193, 32'sd1506,
32'sd747, 32'sd1597, 32'sd682, 32'sd1045, 32'sd878, 32'sd763,
32'sd1023, 32'sd1866, 32'sd1290, 32'sd1979, 32'sd1490, 32'sd1188,
32'sd238, 32'sd1830, 32'sd198, 32'sd724, 32'sd947, 32'sd1294,
32'sd314, 32'sd1480, 32'sd593, 32'sd1809, 32'sd1628, 32'sd508,
32'sd971, 32'sd694, 32'sd1484, 32'sd224, 32'sd662, 32'sd1293,
32'sd967, 32'sd1181, 32'sd674, 32'sd1843, 32'sd977, 32'sd1579,
32'sd820, 32'sd1494, 32'sd238, 32'sd234, 32'sd530, 32'sd979,
32'sd286, 32'sd289, 32'sd295, 32'sd1171, 32'sd817, 32'sd1357,
32'sd922, 32'sd430, 32'sd723, 32'sd1838, 32'sd1172, 32'sd1727,
32'sd146, 32'sd1015, 32'sd1944, 32'sd713, 32'sd536, 32'sd414,
32'sd255, 32'sd1884, 32'sd1353, 32'sd656, 32'sd1656, 32'sd920,
32'sd917, 32'sd1418, 32'sd1637, 32'sd557, 32'sd437, 32'sd1066,
32'sd226, 32'sd1818, 32'sd921, 32'sd762, 32'sd115, 32'sd1885,
32'sd1050, 32'sd472, 32'sd582, 32'sd1882, 32'sd1858, 32'sd1983,
32'sd388, 32'sd1242, 32'sd1202, 32'sd742, 32'sd1582, 32'sd630,
32'sd707, 32'sd1024, 32'sd451, 32'sd1642, 32'sd1342, 32'sd874,
32'sd1962, 32'sd916, 32'sd1356, 32'sd1820, 32'sd1515, 32'sd552,
32'sd1934, 32'sd1177, 32'sd1190, 32'sd1231, 32'sd887, 32'sd1360,
32'sd387, 32'sd998, 32'sd1780, 32'sd356, 32'sd754, 32'sd1614,
32'sd1537, 32'sd134, 32'sd299, 32'sd645, 32'sd887, 32'sd1496,
32'sd1394, 32'sd1168, 32'sd1097, 32'sd543, 32'sd521, 32'sd965,
32'sd1045, 32'sd805, 32'sd1145, 32'sd866, 32'sd1857, 32'sd1195,
32'sd342, 32'sd1374, 32'sd789, 32'sd1519, 32'sd528, 32'sd1365,
32'sd208, 32'sd1553, 32'sd1857, 32'sd475, 32'sd1037, 32'sd1866,
32'sd166, 32'sd686, 32'sd1331, 32'sd1833, 32'sd1764, 32'sd684,
32'sd1460, 32'sd1824, 32'sd1602, 32'sd1578, 32'sd396, 32'sd1103,
32'sd1817, 32'sd1020, 32'sd1858, 32'sd1931, 32'sd757, 32'sd270,
32'sd984, 32'sd594, 32'sd1225, 32'sd1217, 32'sd1517, 32'sd1334,
32'sd1312, 32'sd485, 32'sd369, 32'sd1677, 32'sd290, 32'sd624,
32'sd434, 32'sd171, 32'sd1667, 32'sd1284, 32'sd240, 32'sd952,
32'sd295, 32'sd1647, 32'sd718, 32'sd1962, 32'sd520, 32'sd1641,
32'sd365, 32'sd1387, 32'sd1123, 32'sd847, 32'sd185, 32'sd1522,
32'sd324, 32'sd1954, 32'sd338, 32'sd1011, 32'sd146, 32'sd1980,
32'sd176, 32'sd352, 32'sd997, 32'sd1678, 32'sd551, 32'sd1107,
32'sd324, 32'sd1904, 32'sd1021, 32'sd189, 32'sd1158, 32'sd681,
32'sd690, 32'sd1346, 32'sd787, 32'sd1505, 32'sd1560, 32'sd341,
32'sd1278, 32'sd131, 32'sd475, 32'sd428, 32'sd1851, 32'sd461,
32'sd1020, 32'sd791, 32'sd1318, 32'sd1466, 32'sd1858, 32'sd1327,
32'sd1806, 32'sd1040, 32'sd359, 32'sd400, 32'sd1670, 32'sd1628,
32'sd958, 32'sd503, 32'sd1656, 32'sd833, 32'sd1200, 32'sd848,
32'sd1601, 32'sd1673, 32'sd417, 32'sd480, 32'sd959, 32'sd1970,
32'sd1003, 32'sd729, 32'sd226, 32'sd351, 32'sd1975, 32'sd1797,
32'sd1575, 32'sd634, 32'sd1825, 32'sd312, 32'sd895, 32'sd1807,
32'sd1676, 32'sd273, 32'sd312, 32'sd1258, 32'sd1915, 32'sd1904,
32'sd1286, 32'sd811, 32'sd413, 32'sd874, 32'sd1882, 32'sd1027,
32'sd1502, 32'sd349, 32'sd1296, 32'sd373, 32'sd433, 32'sd779,
32'sd1526, 32'sd1342, 32'sd537, 32'sd1702, 32'sd1870, 32'sd343,
32'sd804, 32'sd459, 32'sd313, 32'sd1499, 32'sd1827, 32'sd968,
32'sd1278, 32'sd824, 32'sd1620, 32'sd1623, 32'sd103, 32'sd386,
32'sd818, 32'sd162, 32'sd972, 32'sd1557, 32'sd1082, 32'sd1709,
32'sd1330, 32'sd912, 32'sd1755, 32'sd984, 32'sd266, 32'sd1650,
32'sd944, 32'sd1851, 32'sd439, 32'sd637, 32'sd798, 32'sd1767,
32'sd937, 32'sd987, 32'sd1845, 32'sd1557, 32'sd1484, 32'sd861,
32'sd246, 32'sd922, 32'sd1576, 32'sd1735, 32'sd916, 32'sd787,
32'sd1215, 32'sd880, 32'sd625, 32'sd922, 32'sd1657, 32'sd169,
32'sd354, 32'sd1656, 32'sd1533, 32'sd1367, 32'sd1905, 32'sd1147,
32'sd107, 32'sd1415, 32'sd1250, 32'sd1054, 32'sd1111, 32'sd148,
32'sd500, 32'sd1424, 32'sd1123, 32'sd1182, 32'sd368, 32'sd103,
32'sd1200, 32'sd1914, 32'sd120, 32'sd634, 32'sd758, 32'sd425,
32'sd1688, 32'sd363, 32'sd1123, 32'sd989, 32'sd1002, 32'sd1045,
32'sd212, 32'sd631, 32'sd1921, 32'sd796, 32'sd171, 32'sd1766,
32'sd141, 32'sd662, 32'sd304, 32'sd920, 32'sd537, 32'sd1299,
32'sd859, 32'sd1273, 32'sd127, 32'sd753, 32'sd1647, 32'sd400,
32'sd481, 32'sd1230, 32'sd1444, 32'sd1861, 32'sd1516, 32'sd361,
32'sd1041, 32'sd1559, 32'sd1563, 32'sd309, 32'sd349, 32'sd129,
32'sd1312, 32'sd1907, 32'sd124, 32'sd1442, 32'sd1007, 32'sd566,
32'sd228, 32'sd647, 32'sd1978, 32'sd1492, 32'sd1519, 32'sd119,
32'sd644, 32'sd1657, 32'sd1662, 32'sd1234, 32'sd1702, 32'sd1628,
32'sd124, 32'sd443, 32'sd1273, 32'sd498, 32'sd994, 32'sd1613,
32'sd1378, 32'sd1656, 32'sd1249, 32'sd1577, 32'sd979, 32'sd1328,
32'sd1103, 32'sd724, 32'sd668, 32'sd1907, 32'sd1066, 32'sd1730,
32'sd1643, 32'sd1056, 32'sd1962, 32'sd831, 32'sd1827, 32'sd1365,
32'sd907, 32'sd1247, 32'sd1539, 32'sd1023, 32'sd1661, 32'sd719,
32'sd1830, 32'sd327, 32'sd1778, 32'sd123, 32'sd319, 32'sd1895,
32'sd141, 32'sd1006, 32'sd293, 32'sd451, 32'sd629, 32'sd794,
32'sd1860, 32'sd1290, 32'sd247, 32'sd1490, 32'sd934, 32'sd1120,
32'sd1444, 32'sd408, 32'sd1786, 32'sd1034, 32'sd1532, 32'sd1737,
32'sd912, 32'sd976, 32'sd788, 32'sd534, 32'sd326, 32'sd1959,
32'sd923, 32'sd232, 32'sd142, 32'sd1444, 32'sd284, 32'sd910,
32'sd1380, 32'sd1484, 32'sd871, 32'sd1420, 32'sd775, 32'sd1606,
32'sd1736, 32'sd1394, 32'sd1582, 32'sd367, 32'sd1611, 32'sd316,
32'sd409, 32'sd1934, 32'sd1511, 32'sd1706, 32'sd767, 32'sd305,
32'sd645, 32'sd1350, 32'sd1765, 32'sd810, 32'sd1010, 32'sd765,
32'sd508, 32'sd1147, 32'sd1864, 32'sd1584, 32'sd772, 32'sd1938,
32'sd1147, 32'sd753, 32'sd163, 32'sd150, 32'sd1207, 32'sd1988,
32'sd1337, 32'sd1497, 32'sd1529, 32'sd1201, 32'sd116, 32'sd1824,
32'sd405, 32'sd1847, 32'sd1212, 32'sd1744, 32'sd817, 32'sd1227,
32'sd1207, 32'sd160, 32'sd1173, 32'sd811, 32'sd562, 32'sd516,
32'sd1628, 32'sd779, 32'sd182, 32'sd1939, 32'sd1608, 32'sd1527,
32'sd1837, 32'sd1531, 32'sd1186, 32'sd1988, 32'sd1098, 32'sd587,
32'sd228, 32'sd1295, 32'sd1366, 32'sd1156, 32'sd600, 32'sd1576,
32'sd1725, 32'sd1462, 32'sd1526, 32'sd1369, 32'sd982, 32'sd1531,
32'sd1081, 32'sd921, 32'sd704, 32'sd1726, 32'sd1645, 32'sd794,
32'sd855, 32'sd1295, 32'sd828, 32'sd1931, 32'sd308, 32'sd345,
32'sd1486, 32'sd1950, 32'sd141, 32'sd1292, 32'sd1887, 32'sd1203,
32'sd341, 32'sd1603, 32'sd1290, 32'sd212, 32'sd854, 32'sd207,
32'sd689, 32'sd1046, 32'sd1267, 32'sd1034, 32'sd827, 32'sd686,
32'sd1776, 32'sd364, 32'sd1568, 32'sd100, 32'sd502, 32'sd124,
32'sd860, 32'sd1269, 32'sd1817, 32'sd999, 32'sd603, 32'sd573,
32'sd416, 32'sd1611, 32'sd123, 32'sd1163, 32'sd1391, 32'sd1724,
32'sd1270, 32'sd734, 32'sd1871, 32'sd162, 32'sd405, 32'sd1903,
32'sd382, 32'sd1889, 32'sd228, 32'sd486, 32'sd823, 32'sd239,
32'sd1160, 32'sd647, 32'sd730, 32'sd1743, 32'sd1458, 32'sd244,
32'sd1203, 32'sd1983, 32'sd1980, 32'sd675, 32'sd132, 32'sd1158,
32'sd924, 32'sd591, 32'sd1496, 32'sd508, 32'sd1257, 32'sd1785,
32'sd1061, 32'sd1680, 32'sd1729, 32'sd872, 32'sd770, 32'sd1919,
32'sd1521, 32'sd1728, 32'sd459, 32'sd790, 32'sd624, 32'sd1481,
32'sd1428, 32'sd1843, 32'sd775, 32'sd1691, 32'sd749, 32'sd525,
32'sd1505, 32'sd1197, 32'sd215, 32'sd1408, 32'sd1444, 32'sd1537,
32'sd682, 32'sd247, 32'sd344, 32'sd627, 32'sd932, 32'sd951,
32'sd270, 32'sd1478, 32'sd223, 32'sd511, 32'sd1147, 32'sd1353,
32'sd1183, 32'sd1877, 32'sd687, 32'sd1283, 32'sd1850, 32'sd1456,
32'sd1706, 32'sd1604, 32'sd681, 32'sd1840, 32'sd1480, 32'sd1180,
32'sd1793, 32'sd158, 32'sd813, 32'sd324, 32'sd925, 32'sd1776,
32'sd1557, 32'sd769, 32'sd1873, 32'sd1455, 32'sd1969, 32'sd1440,
32'sd560, 32'sd339, 32'sd1857, 32'sd1151, 32'sd1753, 32'sd1891,
32'sd1494, 32'sd1235, 32'sd1548, 32'sd334, 32'sd1407, 32'sd710,
32'sd414, 32'sd508, 32'sd521, 32'sd872, 32'sd1435, 32'sd511,
32'sd1821, 32'sd1534, 32'sd610, 32'sd1139, 32'sd596, 32'sd1534,
32'sd1425, 32'sd912, 32'sd1128, 32'sd741, 32'sd1531, 32'sd1120,
32'sd1092, 32'sd853, 32'sd1324, 32'sd1257, 32'sd1875, 32'sd1558,
32'sd627, 32'sd921, 32'sd1213, 32'sd1769, 32'sd1727, 32'sd1470,
32'sd1897, 32'sd117, 32'sd1621, 32'sd275, 32'sd811, 32'sd1695,
32'sd661, 32'sd1226, 32'sd493, 32'sd1338, 32'sd1530, 32'sd918,
32'sd1106, 32'sd273, 32'sd739, 32'sd723, 32'sd1581, 32'sd370,
32'sd641, 32'sd1129, 32'sd1807, 32'sd1000, 32'sd885, 32'sd1823,
32'sd746, 32'sd1016, 32'sd1726, 32'sd659, 32'sd891, 32'sd1018,
32'sd682, 32'sd815, 32'sd171, 32'sd1384, 32'sd156, 32'sd1935,
32'sd800, 32'sd987, 32'sd1585, 32'sd1678, 32'sd260, 32'sd1352,
32'sd1308, 32'sd1434, 32'sd1466, 32'sd1086, 32'sd754, 32'sd949,
32'sd1946, 32'sd1979, 32'sd1182, 32'sd378, 32'sd1035, 32'sd1712,
32'sd1530, 32'sd303, 32'sd1894, 32'sd1081, 32'sd302, 32'sd1920,
32'sd200, 32'sd851, 32'sd439, 32'sd825, 32'sd767, 32'sd1028,
32'sd1123, 32'sd1235, 32'sd1300, 32'sd651, 32'sd752, 32'sd170,
32'sd1284, 32'sd996, 32'sd1628, 32'sd1271, 32'sd1949, 32'sd409,
32'sd1267, 32'sd683, 32'sd1148, 32'sd1574, 32'sd594, 32'sd1938,
32'sd259, 32'sd198, 32'sd1437, 32'sd1885, 32'sd444, 32'sd1512,
32'sd1443, 32'sd1022, 32'sd1431, 32'sd1355, 32'sd1980, 32'sd336,
32'sd754, 32'sd1630, 32'sd422, 32'sd1124, 32'sd456, 32'sd716,
32'sd1511, 32'sd1693, 32'sd1356, 32'sd438, 32'sd1772, 32'sd1408,
32'sd1832, 32'sd315, 32'sd321, 32'sd1554, 32'sd514, 32'sd1134,
32'sd491, 32'sd372, 32'sd419, 32'sd871, 32'sd212, 32'sd627,
32'sd1836, 32'sd671, 32'sd1322, 32'sd1468, 32'sd1029, 32'sd812,
32'sd547, 32'sd701, 32'sd152, 32'sd1431, 32'sd789, 32'sd1482,
32'sd162, 32'sd608, 32'sd814, 32'sd384, 32'sd1595, 32'sd1118,
32'sd678, 32'sd1713, 32'sd1804, 32'sd733, 32'sd986, 32'sd1842,
32'sd440, 32'sd761, 32'sd1470, 32'sd1230, 32'sd1220, 32'sd1744,
32'sd1852, 32'sd1217, 32'sd667, 32'sd826, 32'sd757, 32'sd1437,
32'sd344, 32'sd1940, 32'sd1371, 32'sd1110, 32'sd1323, 32'sd1657,
32'sd1384, 32'sd1851, 32'sd435, 32'sd658, 32'sd767, 32'sd1568,
32'sd413, 32'sd1203, 32'sd730, 32'sd888, 32'sd1463, 32'sd1107,
32'sd1117, 32'sd142, 32'sd1005, 32'sd1056, 32'sd1862, 32'sd1681,
32'sd725, 32'sd1854, 32'sd1118, 32'sd454, 32'sd415, 32'sd849,
32'sd478, 32'sd1324, 32'sd923, 32'sd327, 32'sd1847, 32'sd1940,
32'sd304, 32'sd1938, 32'sd1596, 32'sd895, 32'sd487, 32'sd626,
32'sd1500, 32'sd1278, 32'sd853, 32'sd1945, 32'sd1142, 32'sd1877,
32'sd1165, 32'sd1211, 32'sd989, 32'sd1487, 32'sd1263, 32'sd267,
32'sd877, 32'sd1317, 32'sd113, 32'sd960, 32'sd516, 32'sd1515,
32'sd788, 32'sd191, 32'sd499, 32'sd985, 32'sd1269, 32'sd1581,
32'sd1251, 32'sd654, 32'sd686, 32'sd131, 32'sd861, 32'sd700,
32'sd1071, 32'sd1344, 32'sd1901, 32'sd1452, 32'sd1524, 32'sd1533,
32'sd386, 32'sd301, 32'sd260, 32'sd324, 32'sd400, 32'sd537,
32'sd1957, 32'sd1824, 32'sd1763, 32'sd410, 32'sd1456, 32'sd574,
32'sd195, 32'sd1636, 32'sd1090, 32'sd1434, 32'sd155, 32'sd329,
32'sd1356, 32'sd1401, 32'sd1737, 32'sd594, 32'sd1184, 32'sd1122,
32'sd1613, 32'sd125, 32'sd1417, 32'sd1069, 32'sd748, 32'sd1718,
32'sd748, 32'sd1058, 32'sd1120, 32'sd411, 32'sd1498, 32'sd718,
32'sd633, 32'sd1781, 32'sd878, 32'sd1049, 32'sd989, 32'sd1985,
32'sd1312, 32'sd1366, 32'sd1701, 32'sd1920, 32'sd434, 32'sd1237,
32'sd783, 32'sd956, 32'sd391, 32'sd1410, 32'sd1386, 32'sd599,
32'sd1101, 32'sd969, 32'sd1292, 32'sd1664, 32'sd555, 32'sd1842,
32'sd496, 32'sd439, 32'sd1070, 32'sd405, 32'sd1837, 32'sd1266,
32'sd1158, 32'sd1879, 32'sd1424, 32'sd1408, 32'sd892, 32'sd1755,
32'sd1104, 32'sd1684, 32'sd617, 32'sd550, 32'sd901, 32'sd199,
32'sd1852, 32'sd714, 32'sd1048, 32'sd480, 32'sd1120, 32'sd1813,
32'sd1162, 32'sd540, 32'sd1597, 32'sd226, 32'sd416, 32'sd1519,
32'sd770, 32'sd1477, 32'sd951, 32'sd1440, 32'sd1893, 32'sd341,
32'sd1281, 32'sd312, 32'sd1588, 32'sd579, 32'sd1709, 32'sd1283,
32'sd826, 32'sd996, 32'sd1946, 32'sd1234, 32'sd816, 32'sd1078,
32'sd1792, 32'sd1935, 32'sd1035, 32'sd162, 32'sd1553, 32'sd587,
32'sd928, 32'sd492, 32'sd1373, 32'sd1068, 32'sd719, 32'sd1789,
32'sd1629, 32'sd401, 32'sd329, 32'sd460, 32'sd1444, 32'sd625,
32'sd820, 32'sd777, 32'sd1694, 32'sd805, 32'sd1373, 32'sd992,
32'sd249, 32'sd1821, 32'sd924, 32'sd797, 32'sd164, 32'sd1884,
32'sd1541, 32'sd578, 32'sd883, 32'sd639, 32'sd1898, 32'sd1261,
32'sd1058, 32'sd1946, 32'sd1331, 32'sd1534, 32'sd1130, 32'sd149,
32'sd1975, 32'sd1949, 32'sd1549, 32'sd1153, 32'sd1875, 32'sd155,
32'sd1002, 32'sd878, 32'sd1213, 32'sd698, 32'sd1565, 32'sd589,
32'sd918, 32'sd233, 32'sd901, 32'sd1043, 32'sd507, 32'sd871,
32'sd1531, 32'sd1448, 32'sd1203, 32'sd585, 32'sd1402, 32'sd1103,
32'sd120, 32'sd1764, 32'sd1680, 32'sd1568, 32'sd770, 32'sd566,
32'sd417, 32'sd1515, 32'sd169, 32'sd527, 32'sd588, 32'sd300,
32'sd997, 32'sd1013, 32'sd908, 32'sd1925, 32'sd1488, 32'sd125,
32'sd1550, 32'sd150, 32'sd282, 32'sd551, 32'sd417, 32'sd443,
32'sd1868, 32'sd293, 32'sd219, 32'sd708, 32'sd894, 32'sd447,
32'sd994, 32'sd1566, 32'sd189, 32'sd1086, 32'sd1821, 32'sd1360,
32'sd835, 32'sd650, 32'sd1738, 32'sd348, 32'sd349, 32'sd1328,
32'sd1443, 32'sd1972, 32'sd246, 32'sd1263, 32'sd205, 32'sd567,
32'sd1327, 32'sd1650, 32'sd721, 32'sd776, 32'sd1249, 32'sd1744,
32'sd478, 32'sd624, 32'sd873, 32'sd835, 32'sd177, 32'sd529,
32'sd584, 32'sd178, 32'sd910, 32'sd1629, 32'sd716, 32'sd1431,
32'sd521, 32'sd1498, 32'sd1283, 32'sd1505, 32'sd1665, 32'sd858,
32'sd932, 32'sd1535, 32'sd1937, 32'sd939, 32'sd650, 32'sd1982,
32'sd1776, 32'sd434, 32'sd328, 32'sd547, 32'sd1840, 32'sd835,
32'sd143, 32'sd394, 32'sd526, 32'sd455, 32'sd614, 32'sd1982,
32'sd1866, 32'sd197, 32'sd1034, 32'sd1146, 32'sd183, 32'sd1499,
32'sd249, 32'sd839, 32'sd1229, 32'sd804, 32'sd1865, 32'sd552,
32'sd317, 32'sd965, 32'sd424, 32'sd1537, 32'sd381, 32'sd500,
32'sd1586, 32'sd1702, 32'sd274, 32'sd171, 32'sd1170, 32'sd981,
32'sd440, 32'sd1992, 32'sd623, 32'sd1242, 32'sd412, 32'sd374,
32'sd344, 32'sd1018, 32'sd165, 32'sd1889, 32'sd885, 32'sd1271,
32'sd1318, 32'sd1437, 32'sd344, 32'sd1467, 32'sd966, 32'sd1618,
32'sd1100, 32'sd1039, 32'sd931, 32'sd757, 32'sd361, 32'sd809,
32'sd1721, 32'sd1001, 32'sd1512, 32'sd713, 32'sd836, 32'sd1327,
32'sd1473, 32'sd1327, 32'sd1646, 32'sd746, 32'sd103, 32'sd669,
32'sd1578, 32'sd106, 32'sd1091, 32'sd1188, 32'sd1540, 32'sd1495,
32'sd519, 32'sd1533, 32'sd618, 32'sd1137, 32'sd1829, 32'sd1038,
32'sd1994, 32'sd1379, 32'sd302, 32'sd1451, 32'sd1507, 32'sd1238,
32'sd572, 32'sd1576, 32'sd1406, 32'sd381, 32'sd1308, 32'sd1787,
32'sd1229, 32'sd1480, 32'sd1280, 32'sd833, 32'sd1832, 32'sd1517,
32'sd1625, 32'sd1552, 32'sd244, 32'sd1924, 32'sd1409, 32'sd1707,
32'sd126, 32'sd974, 32'sd1525, 32'sd1622, 32'sd832, 32'sd290,
32'sd928, 32'sd227, 32'sd1619, 32'sd654, 32'sd1215, 32'sd1611,
32'sd605, 32'sd946, 32'sd1774, 32'sd1139, 32'sd183, 32'sd1723,
32'sd901, 32'sd1602, 32'sd1434, 32'sd1645, 32'sd437, 32'sd707,
32'sd512, 32'sd1010, 32'sd821, 32'sd1005, 32'sd112, 32'sd650,
32'sd485, 32'sd1190, 32'sd772, 32'sd1426, 32'sd713, 32'sd1334,
32'sd1110, 32'sd1275, 32'sd316, 32'sd1465, 32'sd1572, 32'sd110,
32'sd471, 32'sd517, 32'sd1387, 32'sd1104, 32'sd510, 32'sd343,
32'sd1657, 32'sd1863, 32'sd525, 32'sd785, 32'sd1951, 32'sd324,
32'sd1911, 32'sd462, 32'sd171, 32'sd1582, 32'sd943, 32'sd951,
32'sd111, 32'sd1424, 32'sd1820, 32'sd1698, 32'sd469, 32'sd1939,
32'sd1947, 32'sd837, 32'sd205, 32'sd645, 32'sd1616, 32'sd1391,
32'sd1999, 32'sd750, 32'sd1091, 32'sd1425, 32'sd1330, 32'sd1336,
32'sd448, 32'sd178, 32'sd1515, 32'sd175, 32'sd540, 32'sd1068,
32'sd533, 32'sd1993, 32'sd1012, 32'sd641, 32'sd1769, 32'sd1274,
32'sd1431, 32'sd1061, 32'sd1874, 32'sd471, 32'sd454, 32'sd421,
32'sd277, 32'sd1827, 32'sd704, 32'sd278, 32'sd1327, 32'sd967,
32'sd221, 32'sd355, 32'sd1529, 32'sd663, 32'sd144, 32'sd158,
32'sd589, 32'sd823, 32'sd1489, 32'sd1152, 32'sd103, 32'sd1292,
32'sd1319, 32'sd1982, 32'sd597, 32'sd1051, 32'sd728, 32'sd534,
32'sd1718, 32'sd965, 32'sd432, 32'sd549, 32'sd1252, 32'sd1868,
32'sd112, 32'sd1010, 32'sd931, 32'sd1785, 32'sd170, 32'sd523,
32'sd848, 32'sd1854, 32'sd826, 32'sd893, 32'sd1999, 32'sd1311,
32'sd424, 32'sd773, 32'sd1941, 32'sd1509, 32'sd1247, 32'sd1589,
32'sd916, 32'sd1553, 32'sd250, 32'sd713, 32'sd1445, 32'sd1532,
32'sd774, 32'sd1695, 32'sd1139, 32'sd772, 32'sd1547, 32'sd735,
32'sd1940, 32'sd1479, 32'sd1339, 32'sd1689, 32'sd375, 32'sd1837,
32'sd1287, 32'sd553, 32'sd1999, 32'sd156, 32'sd948, 32'sd800,
32'sd1731, 32'sd586, 32'sd330, 32'sd728, 32'sd1551, 32'sd1348,
32'sd965, 32'sd1497, 32'sd550, 32'sd1759, 32'sd1152, 32'sd614,
32'sd1488, 32'sd155, 32'sd1724, 32'sd339, 32'sd1511, 32'sd1352,
32'sd360, 32'sd1838, 32'sd1966, 32'sd1036, 32'sd271, 32'sd139,
32'sd190, 32'sd1060, 32'sd463, 32'sd292, 32'sd1149, 32'sd1757,
32'sd585, 32'sd444, 32'sd339, 32'sd441, 32'sd1577, 32'sd1296,
32'sd750, 32'sd214, 32'sd1382, 32'sd1986, 32'sd1303, 32'sd1116,
32'sd1243, 32'sd451, 32'sd1095, 32'sd1929, 32'sd342, 32'sd691,
32'sd1769, 32'sd1301, 32'sd1390, 32'sd1303, 32'sd296, 32'sd1928,
32'sd1845, 32'sd1844, 32'sd1344, 32'sd744, 32'sd1706, 32'sd638,
32'sd1555, 32'sd651, 32'sd835, 32'sd1025, 32'sd1182, 32'sd838,
32'sd532, 32'sd233, 32'sd339, 32'sd852, 32'sd1987, 32'sd648,
32'sd1511, 32'sd740, 32'sd310, 32'sd435, 32'sd1111, 32'sd1803,
32'sd301, 32'sd1366, 32'sd1312, 32'sd363, 32'sd1463, 32'sd454,
32'sd1173, 32'sd720, 32'sd1052, 32'sd928, 32'sd1138, 32'sd774,
32'sd160, 32'sd1460, 32'sd1629, 32'sd729, 32'sd898, 32'sd387,
32'sd1208, 32'sd1713, 32'sd1320, 32'sd1245, 32'sd1723, 32'sd1791,
32'sd1930, 32'sd1893, 32'sd529, 32'sd1591, 32'sd1407, 32'sd768,
32'sd1399, 32'sd1676, 32'sd1740, 32'sd431, 32'sd689, 32'sd1566,
32'sd1789, 32'sd661, 32'sd149, 32'sd1034, 32'sd321, 32'sd421,
32'sd181, 32'sd206, 32'sd883, 32'sd910, 32'sd1608, 32'sd1476,
32'sd1164, 32'sd1903, 32'sd1445, 32'sd767, 32'sd1835, 32'sd626,
32'sd1047, 32'sd1132, 32'sd489, 32'sd923, 32'sd1700, 32'sd981,
32'sd1138, 32'sd116, 32'sd405, 32'sd913, 32'sd1213, 32'sd1970,
32'sd1807, 32'sd1785, 32'sd620, 32'sd502, 32'sd1024, 32'sd674,
32'sd960, 32'sd1032, 32'sd1066, 32'sd816, 32'sd386, 32'sd468,
32'sd1006, 32'sd472, 32'sd1317, 32'sd624, 32'sd458, 32'sd826,
32'sd769, 32'sd1619, 32'sd196, 32'sd1323, 32'sd1451, 32'sd1667,
32'sd763, 32'sd506, 32'sd443, 32'sd831, 32'sd136, 32'sd1270,
32'sd1205, 32'sd552, 32'sd760, 32'sd1904, 32'sd415, 32'sd924,
32'sd500, 32'sd349, 32'sd101, 32'sd1185, 32'sd1476, 32'sd1670,
32'sd1071, 32'sd834, 32'sd130, 32'sd199, 32'sd1641, 32'sd506,
32'sd1234, 32'sd1495, 32'sd923, 32'sd1196, 32'sd1774, 32'sd1184,
32'sd1462, 32'sd1025, 32'sd1793, 32'sd1779, 32'sd1966, 32'sd428,
32'sd412, 32'sd988, 32'sd330, 32'sd239, 32'sd1363, 32'sd887,
32'sd577, 32'sd598, 32'sd1938, 32'sd234, 32'sd679, 32'sd639,
32'sd1957, 32'sd1897, 32'sd1952, 32'sd263, 32'sd956, 32'sd292,
32'sd731, 32'sd934, 32'sd1929, 32'sd266, 32'sd1263, 32'sd944,
32'sd1350, 32'sd1241, 32'sd1173, 32'sd312, 32'sd1125, 32'sd1427,
32'sd944, 32'sd1394, 32'sd1856, 32'sd1402, 32'sd305, 32'sd1554,
32'sd375, 32'sd1545, 32'sd1915, 32'sd306, 32'sd620, 32'sd122,
32'sd1714, 32'sd1198, 32'sd1010, 32'sd1121, 32'sd1442, 32'sd1902,
32'sd1612, 32'sd893, 32'sd668, 32'sd556, 32'sd414, 32'sd1002,
32'sd866, 32'sd375, 32'sd1496, 32'sd1305, 32'sd557, 32'sd1899,
32'sd1885, 32'sd1970, 32'sd1176, 32'sd631, 32'sd1284, 32'sd1157,
32'sd1441, 32'sd449, 32'sd1101, 32'sd1265, 32'sd557, 32'sd1494,
32'sd933, 32'sd1867, 32'sd1302, 32'sd104, 32'sd965, 32'sd763,
32'sd658, 32'sd1700, 32'sd1896, 32'sd1668, 32'sd1891, 32'sd1196,
32'sd774, 32'sd289, 32'sd1078, 32'sd518, 32'sd1039, 32'sd1750,
32'sd1281, 32'sd897, 32'sd838, 32'sd1459, 32'sd1955, 32'sd973,
32'sd1105, 32'sd485, 32'sd695, 32'sd1935, 32'sd778, 32'sd1480,
32'sd1146, 32'sd1361, 32'sd901, 32'sd217, 32'sd1913, 32'sd971,
32'sd1901, 32'sd1159, 32'sd1619, 32'sd259, 32'sd1198, 32'sd1578,
32'sd1221, 32'sd144, 32'sd758, 32'sd1486, 32'sd1126, 32'sd595,
32'sd1720, 32'sd1091, 32'sd107, 32'sd929, 32'sd316, 32'sd494,
32'sd1086, 32'sd1155, 32'sd1080, 32'sd238, 32'sd1914, 32'sd806,
32'sd723, 32'sd1764, 32'sd943, 32'sd427, 32'sd1890, 32'sd702,
32'sd708, 32'sd419, 32'sd1944, 32'sd1237, 32'sd873, 32'sd1638,
32'sd1821, 32'sd1089, 32'sd1264, 32'sd181, 32'sd1990, 32'sd954,
32'sd864, 32'sd569, 32'sd1984, 32'sd843, 32'sd299, 32'sd1576,
32'sd942, 32'sd1316, 32'sd1852, 32'sd1483, 32'sd1069, 32'sd401,
32'sd1071, 32'sd1245, 32'sd1947, 32'sd639, 32'sd430, 32'sd1368,
32'sd1465, 32'sd697, 32'sd534, 32'sd1675, 32'sd1506, 32'sd1342,
32'sd1667, 32'sd1595, 32'sd938, 32'sd895, 32'sd881, 32'sd372,
32'sd967, 32'sd152, 32'sd415, 32'sd692, 32'sd335, 32'sd1955,
32'sd1233, 32'sd585, 32'sd581, 32'sd389, 32'sd1795, 32'sd1367,
32'sd1161, 32'sd278, 32'sd401, 32'sd424, 32'sd1115, 32'sd1820,
32'sd652, 32'sd468, 32'sd1197, 32'sd1772, 32'sd381, 32'sd1821,
32'sd829, 32'sd1280, 32'sd345, 32'sd1865, 32'sd922, 32'sd881,
32'sd1171, 32'sd324, 32'sd1489, 32'sd984, 32'sd773, 32'sd798,
32'sd980, 32'sd463, 32'sd1790, 32'sd1962, 32'sd888, 32'sd545,
32'sd1908, 32'sd1276, 32'sd1433, 32'sd150, 32'sd398, 32'sd713,
32'sd1499, 32'sd539, 32'sd996, 32'sd571, 32'sd1238, 32'sd1355,
32'sd1836, 32'sd520, 32'sd132, 32'sd215, 32'sd1272, 32'sd266,
32'sd1276, 32'sd483, 32'sd880, 32'sd1729, 32'sd1137, 32'sd1797,
32'sd394, 32'sd1664, 32'sd186, 32'sd1809, 32'sd219, 32'sd1498,
32'sd734, 32'sd1222, 32'sd1941, 32'sd812, 32'sd270, 32'sd1335,
32'sd520, 32'sd1610, 32'sd887, 32'sd1705, 32'sd1371, 32'sd1391,
32'sd1830, 32'sd1649, 32'sd1941, 32'sd1942, 32'sd433, 32'sd466,
32'sd221, 32'sd1576, 32'sd1066, 32'sd356, 32'sd1973, 32'sd1957,
32'sd821, 32'sd599, 32'sd304, 32'sd884, 32'sd1326, 32'sd1119,
32'sd1493, 32'sd1317, 32'sd1290, 32'sd1010, 32'sd701, 32'sd1601,
32'sd1607, 32'sd991, 32'sd1931, 32'sd858, 32'sd146, 32'sd1518,
32'sd1490, 32'sd1614, 32'sd1755, 32'sd1504, 32'sd174, 32'sd359,
32'sd1915, 32'sd681, 32'sd499, 32'sd1341, 32'sd748, 32'sd1959,
32'sd522, 32'sd1399, 32'sd149, 32'sd1893, 32'sd1681, 32'sd246,
32'sd145, 32'sd1126, 32'sd915, 32'sd1098, 32'sd1131, 32'sd1645,
32'sd1212, 32'sd1144, 32'sd999, 32'sd1517, 32'sd1126, 32'sd651,
32'sd277, 32'sd1252, 32'sd1297, 32'sd811, 32'sd1169, 32'sd1910,
32'sd1555, 32'sd412, 32'sd1238, 32'sd1037, 32'sd1970, 32'sd552,
32'sd646, 32'sd1351, 32'sd1682, 32'sd538, 32'sd1771, 32'sd687,
32'sd1762, 32'sd197, 32'sd775, 32'sd1579, 32'sd1379, 32'sd1082,
32'sd1413, 32'sd186, 32'sd1278, 32'sd193, 32'sd1744, 32'sd570,
32'sd1145, 32'sd1634, 32'sd457, 32'sd495, 32'sd1026, 32'sd1264,
32'sd667, 32'sd197, 32'sd1853, 32'sd709, 32'sd564, 32'sd789,
32'sd1591, 32'sd1126, 32'sd809, 32'sd905, 32'sd835, 32'sd670,
32'sd1162, 32'sd1672, 32'sd1745, 32'sd507, 32'sd912, 32'sd1503,
32'sd1499, 32'sd1836, 32'sd891, 32'sd747, 32'sd435, 32'sd1893,
32'sd841, 32'sd1313, 32'sd936, 32'sd901, 32'sd1035, 32'sd673,
32'sd1087, 32'sd130, 32'sd1401, 32'sd315, 32'sd1978, 32'sd1359,
32'sd1494, 32'sd1486, 32'sd1133, 32'sd630, 32'sd758, 32'sd601,
32'sd646, 32'sd417, 32'sd501, 32'sd305, 32'sd1338, 32'sd1838,
32'sd230, 32'sd1143, 32'sd1447, 32'sd573, 32'sd486, 32'sd1532,
32'sd1265, 32'sd634, 32'sd1902, 32'sd1385, 32'sd179, 32'sd423,
32'sd1414, 32'sd434, 32'sd873, 32'sd1398, 32'sd1926, 32'sd129,
32'sd971, 32'sd1795, 32'sd1138, 32'sd376, 32'sd1199, 32'sd1036,
32'sd1582, 32'sd811, 32'sd430, 32'sd1141, 32'sd1095, 32'sd1874,
32'sd740, 32'sd310, 32'sd454, 32'sd1526, 32'sd619, 32'sd1185,
32'sd1683, 32'sd1337, 32'sd1239, 32'sd832, 32'sd587, 32'sd1956,
32'sd1437, 32'sd1052, 32'sd1851, 32'sd566, 32'sd1674, 32'sd311,
32'sd172, 32'sd1510, 32'sd1741, 32'sd1144, 32'sd813, 32'sd1508,
32'sd721, 32'sd1113, 32'sd630, 32'sd1800, 32'sd799, 32'sd762,
32'sd923, 32'sd842, 32'sd751, 32'sd1420, 32'sd1588, 32'sd105,
32'sd1573, 32'sd1925, 32'sd473, 32'sd1464, 32'sd1619, 32'sd758,
32'sd1695, 32'sd1473, 32'sd775, 32'sd131, 32'sd1230, 32'sd1724,
32'sd155, 32'sd1576, 32'sd799, 32'sd1658, 32'sd728, 32'sd962,
32'sd1569, 32'sd1958, 32'sd1055, 32'sd177, 32'sd1601, 32'sd1210,
32'sd1544, 32'sd1595, 32'sd984, 32'sd747, 32'sd1948, 32'sd917,
32'sd1858, 32'sd756, 32'sd911, 32'sd524, 32'sd178, 32'sd125,
32'sd1604, 32'sd1823, 32'sd690, 32'sd338, 32'sd430, 32'sd1729,
32'sd1151, 32'sd1140, 32'sd273, 32'sd127, 32'sd767, 32'sd1788,
32'sd1423, 32'sd1067, 32'sd828, 32'sd1989, 32'sd1501, 32'sd226,
32'sd1972, 32'sd418, 32'sd969, 32'sd1901, 32'sd1514, 32'sd603,
32'sd1861, 32'sd1861, 32'sd1894, 32'sd1164, 32'sd1497, 32'sd877,
32'sd654, 32'sd1880, 32'sd611, 32'sd115, 32'sd919, 32'sd1825,
32'sd1953, 32'sd1906, 32'sd261, 32'sd1472, 32'sd657, 32'sd1822,
32'sd250, 32'sd1670, 32'sd1753, 32'sd919, 32'sd1732, 32'sd1632,
32'sd1604, 32'sd847, 32'sd1807, 32'sd602, 32'sd934, 32'sd1192,
32'sd481, 32'sd698, 32'sd1608, 32'sd1875, 32'sd1316, 32'sd1276,
32'sd1631, 32'sd540, 32'sd1113, 32'sd1233, 32'sd1247, 32'sd1169,
32'sd479, 32'sd609, 32'sd279, 32'sd864, 32'sd148, 32'sd595,
32'sd674, 32'sd554, 32'sd272, 32'sd1717, 32'sd1139, 32'sd1235,
32'sd498, 32'sd1752, 32'sd1089, 32'sd1704, 32'sd685, 32'sd1499,
32'sd967, 32'sd1258, 32'sd720, 32'sd1752, 32'sd443, 32'sd1304,
32'sd1255, 32'sd1583, 32'sd234, 32'sd1982, 32'sd1463, 32'sd1544,
32'sd1545, 32'sd1841, 32'sd1465, 32'sd1495, 32'sd1467, 32'sd1176,
32'sd362, 32'sd1709, 32'sd1690, 32'sd770, 32'sd246, 32'sd141,
32'sd1702, 32'sd606, 32'sd323, 32'sd1756, 32'sd663, 32'sd556,
32'sd125, 32'sd903, 32'sd675, 32'sd547, 32'sd409, 32'sd1446,
32'sd1905, 32'sd794, 32'sd1244, 32'sd606, 32'sd171, 32'sd1999,
32'sd716, 32'sd574, 32'sd665, 32'sd1089, 32'sd873, 32'sd1917,
32'sd1376, 32'sd423, 32'sd1705, 32'sd1937, 32'sd1227, 32'sd1370,
32'sd734, 32'sd1887, 32'sd452, 32'sd1299, 32'sd1198, 32'sd594,
32'sd1541, 32'sd263, 32'sd914, 32'sd1817, 32'sd286, 32'sd105,
32'sd581, 32'sd955, 32'sd1857, 32'sd1507, 32'sd1987, 32'sd290,
32'sd1191, 32'sd187, 32'sd1484, 32'sd1813, 32'sd1450, 32'sd1745,
32'sd1693, 32'sd1894, 32'sd1338, 32'sd1973, 32'sd743, 32'sd144,
32'sd1861, 32'sd658, 32'sd178, 32'sd1219, 32'sd747, 32'sd154,
32'sd1621, 32'sd1240, 32'sd412, 32'sd1460, 32'sd1437, 32'sd1355,
32'sd1349, 32'sd559, 32'sd1317, 32'sd473, 32'sd1199, 32'sd1931,
32'sd374, 32'sd853, 32'sd305, 32'sd1718, 32'sd1562, 32'sd1446,
32'sd1222, 32'sd883, 32'sd866, 32'sd1100, 32'sd1329, 32'sd719,
32'sd853, 32'sd224, 32'sd1637, 32'sd1135, 32'sd1263, 32'sd1892,
32'sd1266, 32'sd1012, 32'sd452, 32'sd1287, 32'sd928, 32'sd1949,
32'sd405, 32'sd568, 32'sd1950, 32'sd847, 32'sd415, 32'sd668,
32'sd443, 32'sd359, 32'sd1087, 32'sd657, 32'sd760, 32'sd1377,
32'sd1847, 32'sd1505, 32'sd1099, 32'sd1269, 32'sd150, 32'sd139,
32'sd808, 32'sd891, 32'sd1058, 32'sd762, 32'sd633, 32'sd314,
32'sd1539, 32'sd1471, 32'sd745, 32'sd797, 32'sd965, 32'sd1755,
32'sd1012, 32'sd1738, 32'sd1835, 32'sd601, 32'sd1272, 32'sd1136,
32'sd1015, 32'sd519, 32'sd1772, 32'sd321, 32'sd1790, 32'sd1757,
32'sd1283, 32'sd969, 32'sd1366, 32'sd1481, 32'sd226, 32'sd777,
32'sd1111, 32'sd1686, 32'sd1678, 32'sd614, 32'sd1370, 32'sd1650,
32'sd118, 32'sd753, 32'sd463, 32'sd1493, 32'sd1748, 32'sd168,
32'sd1642, 32'sd639, 32'sd234, 32'sd1150, 32'sd866, 32'sd1886,
32'sd249, 32'sd661, 32'sd1750, 32'sd1725, 32'sd1857, 32'sd951,
32'sd1067, 32'sd1765, 32'sd1988, 32'sd1306, 32'sd1859, 32'sd758,
32'sd961, 32'sd522, 32'sd1334, 32'sd1906, 32'sd445, 32'sd1132,
32'sd911, 32'sd1468, 32'sd790, 32'sd1312, 32'sd664, 32'sd431,
32'sd1326, 32'sd726, 32'sd203, 32'sd745, 32'sd220, 32'sd429,
32'sd152, 32'sd1024, 32'sd303, 32'sd1409, 32'sd1514, 32'sd491,
32'sd1225, 32'sd779, 32'sd207, 32'sd1231, 32'sd1011, 32'sd925,
32'sd1033, 32'sd1999, 32'sd508, 32'sd634, 32'sd163, 32'sd1556,
32'sd1573, 32'sd776, 32'sd1958, 32'sd886, 32'sd1925, 32'sd1005,
32'sd1338, 32'sd708, 32'sd1168, 32'sd1828, 32'sd1345, 32'sd1048,
32'sd1825, 32'sd1440, 32'sd1072, 32'sd1610, 32'sd1648, 32'sd1832,
32'sd1119, 32'sd1881, 32'sd543, 32'sd1580, 32'sd781, 32'sd362,
32'sd1198, 32'sd1430, 32'sd1588, 32'sd1618, 32'sd924, 32'sd192,
32'sd774, 32'sd1953, 32'sd320, 32'sd1141, 32'sd1221, 32'sd1699,
32'sd640, 32'sd613, 32'sd504, 32'sd139, 32'sd1407, 32'sd1259,
32'sd1790, 32'sd1766, 32'sd1021, 32'sd675, 32'sd1899, 32'sd370,
32'sd966, 32'sd1448, 32'sd688, 32'sd1523, 32'sd937, 32'sd1083,
32'sd747, 32'sd402, 32'sd499, 32'sd427, 32'sd308, 32'sd206,
32'sd1689, 32'sd805, 32'sd983, 32'sd826, 32'sd143, 32'sd884,
32'sd1113, 32'sd1609, 32'sd320, 32'sd592, 32'sd1017, 32'sd743,
32'sd818, 32'sd1319, 32'sd1568, 32'sd1639, 32'sd690, 32'sd1459,
32'sd501, 32'sd1489, 32'sd1200, 32'sd1782, 32'sd169, 32'sd799,
32'sd187, 32'sd495, 32'sd1872, 32'sd1771, 32'sd286, 32'sd394,
32'sd1948, 32'sd1264, 32'sd1495, 32'sd1060, 32'sd1607, 32'sd1312,
32'sd1540, 32'sd811, 32'sd272, 32'sd101, 32'sd1219, 32'sd1723,
32'sd844, 32'sd548, 32'sd714, 32'sd1791, 32'sd1707, 32'sd1797,
32'sd1595, 32'sd264, 32'sd921, 32'sd1432, 32'sd1480, 32'sd1731,
32'sd1616, 32'sd160, 32'sd861, 32'sd1259, 32'sd479, 32'sd1059,
32'sd505, 32'sd1264, 32'sd1402, 32'sd590, 32'sd1583, 32'sd1835,
32'sd1080, 32'sd1436, 32'sd1706, 32'sd664, 32'sd1531, 32'sd167,
32'sd664, 32'sd426, 32'sd920, 32'sd1467, 32'sd158, 32'sd1566,
32'sd624, 32'sd1092, 32'sd446, 32'sd1011, 32'sd524, 32'sd256,
32'sd1326, 32'sd509, 32'sd617, 32'sd718, 32'sd1599, 32'sd1560,
32'sd1288, 32'sd1317, 32'sd180, 32'sd257, 32'sd1291, 32'sd1586,
32'sd100, 32'sd1090, 32'sd563, 32'sd1457, 32'sd296, 32'sd416,
32'sd1520, 32'sd972, 32'sd1663, 32'sd1166, 32'sd763, 32'sd329,
32'sd1507, 32'sd1433, 32'sd1598, 32'sd1907, 32'sd110, 32'sd1527,
32'sd1675, 32'sd246, 32'sd880, 32'sd1568, 32'sd203, 32'sd753,
32'sd874, 32'sd1004, 32'sd1461, 32'sd1743, 32'sd1123, 32'sd1374,
32'sd1875, 32'sd1986, 32'sd420, 32'sd420, 32'sd1474, 32'sd1498,
32'sd1092, 32'sd1541, 32'sd1472, 32'sd1377, 32'sd743, 32'sd1067,
32'sd1227, 32'sd1119, 32'sd1208, 32'sd1578, 32'sd1460, 32'sd945,
32'sd1227, 32'sd237, 32'sd671, 32'sd182, 32'sd1005, 32'sd1321,
32'sd1793, 32'sd1632, 32'sd1834, 32'sd545, 32'sd484, 32'sd784,
32'sd1023, 32'sd107, 32'sd473, 32'sd1651, 32'sd1584, 32'sd1592,
32'sd1548, 32'sd1218, 32'sd1127, 32'sd1644, 32'sd696, 32'sd1410,
32'sd1282, 32'sd1992, 32'sd1941, 32'sd509, 32'sd1234, 32'sd1509,
32'sd284, 32'sd817, 32'sd1851, 32'sd458, 32'sd958, 32'sd1110,
32'sd684, 32'sd1316, 32'sd1268, 32'sd1521, 32'sd1496, 32'sd1697,
32'sd448, 32'sd1877, 32'sd409, 32'sd1110, 32'sd867, 32'sd1200,
32'sd1783, 32'sd1511, 32'sd232, 32'sd409, 32'sd1267, 32'sd796,
32'sd1487, 32'sd586, 32'sd1287, 32'sd1233, 32'sd1590, 32'sd1967,
32'sd665, 32'sd1505, 32'sd1132, 32'sd904, 32'sd1361, 32'sd674,
32'sd106, 32'sd357, 32'sd1511, 32'sd1728, 32'sd1189, 32'sd372,
32'sd961, 32'sd1545, 32'sd568, 32'sd982, 32'sd955, 32'sd1459,
32'sd1014, 32'sd866, 32'sd614, 32'sd931, 32'sd132, 32'sd852,
32'sd1027, 32'sd1990, 32'sd848, 32'sd462, 32'sd1828, 32'sd1848,
32'sd796, 32'sd429, 32'sd460, 32'sd1174, 32'sd1481, 32'sd806,
32'sd558, 32'sd1632, 32'sd955, 32'sd775, 32'sd1871, 32'sd1247,
32'sd763, 32'sd1988, 32'sd523, 32'sd1407, 32'sd456, 32'sd571,
32'sd203, 32'sd432, 32'sd1899, 32'sd1639, 32'sd1222, 32'sd404,
32'sd1463, 32'sd1242, 32'sd1299, 32'sd291, 32'sd171, 32'sd979,
32'sd833, 32'sd1408, 32'sd410, 32'sd1565, 32'sd288, 32'sd572,
32'sd1156, 32'sd286, 32'sd355, 32'sd1960, 32'sd902, 32'sd1395,
32'sd275, 32'sd512, 32'sd1483, 32'sd897, 32'sd500, 32'sd977,
32'sd318, 32'sd278, 32'sd1372, 32'sd1957, 32'sd1939, 32'sd1468,
32'sd465, 32'sd279, 32'sd267, 32'sd894, 32'sd1397, 32'sd1296,
32'sd1667, 32'sd1526, 32'sd417, 32'sd1733, 32'sd1044, 32'sd783,
32'sd1178, 32'sd1932, 32'sd1878, 32'sd997, 32'sd939, 32'sd512,
32'sd134, 32'sd1103, 32'sd433, 32'sd1099, 32'sd185, 32'sd1120,
32'sd477, 32'sd1252, 32'sd884, 32'sd1928, 32'sd808, 32'sd458,
32'sd957, 32'sd695, 32'sd176, 32'sd990, 32'sd356, 32'sd589,
32'sd1419, 32'sd1232, 32'sd434, 32'sd1833, 32'sd1923, 32'sd429,
32'sd950, 32'sd198, 32'sd312, 32'sd1935, 32'sd536, 32'sd1294,
32'sd294, 32'sd1549, 32'sd1248, 32'sd1829, 32'sd1833, 32'sd117,
32'sd1974, 32'sd570, 32'sd1191, 32'sd1042, 32'sd847, 32'sd808,
32'sd703, 32'sd425, 32'sd1952, 32'sd1905, 32'sd715, 32'sd821,
32'sd1991, 32'sd1301, 32'sd1961, 32'sd1407, 32'sd1836, 32'sd1339,
32'sd1394, 32'sd1211, 32'sd1576, 32'sd878, 32'sd444, 32'sd876,
32'sd633, 32'sd1641, 32'sd1289, 32'sd970, 32'sd1831, 32'sd554,
32'sd1956, 32'sd437, 32'sd291, 32'sd1354, 32'sd145, 32'sd363,
32'sd803, 32'sd936, 32'sd1467, 32'sd208, 32'sd379, 32'sd1887,
32'sd1127, 32'sd680, 32'sd1168, 32'sd1325, 32'sd1651, 32'sd756,
32'sd570, 32'sd1233, 32'sd792, 32'sd1625, 32'sd293, 32'sd1899,
32'sd856, 32'sd1903, 32'sd1370, 32'sd1134, 32'sd1696, 32'sd168,
32'sd1551, 32'sd1683, 32'sd817, 32'sd1068, 32'sd1645, 32'sd924,
32'sd1781, 32'sd689, 32'sd1852, 32'sd1924, 32'sd1318, 32'sd1810,
32'sd1101, 32'sd1624, 32'sd583, 32'sd770, 32'sd265, 32'sd1091,
32'sd1163, 32'sd1175, 32'sd1787, 32'sd612, 32'sd944, 32'sd291,
32'sd505, 32'sd845, 32'sd1715, 32'sd1990, 32'sd202, 32'sd1932,
32'sd1312, 32'sd1458, 32'sd989, 32'sd1862, 32'sd602, 32'sd684,
32'sd1193, 32'sd697, 32'sd1858, 32'sd1907, 32'sd850, 32'sd372,
32'sd941, 32'sd1622, 32'sd1085, 32'sd125, 32'sd335, 32'sd1817,
32'sd1469, 32'sd1883, 32'sd551, 32'sd128, 32'sd1657, 32'sd1674,
32'sd1349, 32'sd868, 32'sd1062, 32'sd255, 32'sd662, 32'sd535,
32'sd1253, 32'sd1163, 32'sd1388, 32'sd1296, 32'sd1483, 32'sd362,
32'sd1407, 32'sd804, 32'sd776, 32'sd1174, 32'sd1839, 32'sd337,
32'sd1876, 32'sd948, 32'sd1063, 32'sd580, 32'sd145, 32'sd552,
32'sd1056, 32'sd1715, 32'sd1334, 32'sd447, 32'sd213, 32'sd1222,
32'sd545, 32'sd829, 32'sd228, 32'sd596, 32'sd536, 32'sd490,
32'sd359, 32'sd1717, 32'sd809, 32'sd280, 32'sd850, 32'sd1952,
32'sd1484, 32'sd1155, 32'sd1915, 32'sd404, 32'sd439, 32'sd1026,
32'sd1577, 32'sd1957, 32'sd101, 32'sd499, 32'sd1438, 32'sd1550,
32'sd1014, 32'sd1506, 32'sd1603, 32'sd1060, 32'sd884, 32'sd912,
32'sd963, 32'sd1834, 32'sd1449, 32'sd385, 32'sd1645, 32'sd341,
32'sd1329, 32'sd1748, 32'sd153, 32'sd123, 32'sd1046, 32'sd1352,
32'sd1476, 32'sd221, 32'sd1875, 32'sd1659, 32'sd535, 32'sd249,
32'sd1568, 32'sd1959, 32'sd1047, 32'sd1180, 32'sd1125, 32'sd369,
32'sd317, 32'sd1876, 32'sd1051, 32'sd1710, 32'sd433, 32'sd1235,
32'sd1306, 32'sd125, 32'sd453, 32'sd527, 32'sd556, 32'sd1459,
32'sd1729, 32'sd1912, 32'sd1407, 32'sd355, 32'sd854, 32'sd1317,
32'sd160, 32'sd574, 32'sd804, 32'sd640, 32'sd663, 32'sd1030,
32'sd719, 32'sd721, 32'sd1043, 32'sd711, 32'sd476, 32'sd1776,
32'sd1043, 32'sd1146, 32'sd1809, 32'sd1518, 32'sd788, 32'sd460,
32'sd1324, 32'sd325, 32'sd1719, 32'sd167, 32'sd1838, 32'sd1969,
32'sd476, 32'sd602, 32'sd584, 32'sd858, 32'sd334, 32'sd1088,
32'sd628, 32'sd1586, 32'sd328, 32'sd1740, 32'sd113, 32'sd716,
32'sd716, 32'sd1083, 32'sd1978, 32'sd788, 32'sd1007, 32'sd675,
32'sd372, 32'sd141, 32'sd483, 32'sd1817, 32'sd545, 32'sd940,
32'sd976, 32'sd1328, 32'sd1654, 32'sd1173, 32'sd1588, 32'sd554,
32'sd1831, 32'sd809, 32'sd1219, 32'sd646, 32'sd1509, 32'sd183,
32'sd1335, 32'sd509, 32'sd1948, 32'sd1094, 32'sd647, 32'sd1358,
32'sd491, 32'sd1952, 32'sd1372, 32'sd1398, 32'sd1585, 32'sd1998,
32'sd1110, 32'sd1854, 32'sd1211, 32'sd1174, 32'sd1330, 32'sd1246,
32'sd887, 32'sd1677, 32'sd1134, 32'sd329, 32'sd307, 32'sd1641,
32'sd1598, 32'sd1727, 32'sd577, 32'sd951, 32'sd185, 32'sd1479,
32'sd741, 32'sd545, 32'sd1659, 32'sd852, 32'sd280, 32'sd1816,
32'sd733, 32'sd1894, 32'sd551, 32'sd1819, 32'sd1567, 32'sd1685,
32'sd184, 32'sd1795, 32'sd851, 32'sd1257, 32'sd1545, 32'sd847,
32'sd1823, 32'sd166, 32'sd1770, 32'sd138, 32'sd859, 32'sd1830,
32'sd1907, 32'sd1643, 32'sd1968, 32'sd768, 32'sd808, 32'sd524,
32'sd536, 32'sd417, 32'sd987, 32'sd622, 32'sd1836, 32'sd1060,
32'sd298, 32'sd1787, 32'sd339, 32'sd593, 32'sd1195, 32'sd1855,
32'sd1751, 32'sd397, 32'sd390, 32'sd1724, 32'sd1134, 32'sd1616,
32'sd235, 32'sd999, 32'sd1233, 32'sd475, 32'sd452, 32'sd849,
32'sd387, 32'sd643, 32'sd1817, 32'sd1476, 32'sd1595, 32'sd270,
32'sd1010, 32'sd1731, 32'sd496, 32'sd1745, 32'sd855, 32'sd1781,
32'sd1321, 32'sd1108, 32'sd879, 32'sd1129, 32'sd1686, 32'sd1844,
32'sd1978, 32'sd621, 32'sd1662, 32'sd367, 32'sd1317, 32'sd707,
32'sd689, 32'sd424, 32'sd1326, 32'sd437, 32'sd448, 32'sd217,
32'sd143, 32'sd459, 32'sd1522, 32'sd1462, 32'sd1336, 32'sd722,
32'sd541, 32'sd250, 32'sd616, 32'sd1474, 32'sd780, 32'sd1789,
32'sd753, 32'sd658, 32'sd1752, 32'sd974, 32'sd1428, 32'sd932,
32'sd1825, 32'sd1310, 32'sd802, 32'sd913, 32'sd340, 32'sd1314,
32'sd1027, 32'sd836, 32'sd1738, 32'sd1889, 32'sd1587, 32'sd1852,
32'sd1830, 32'sd772, 32'sd1071, 32'sd841, 32'sd205, 32'sd1446,
32'sd1764, 32'sd1020, 32'sd621, 32'sd1497, 32'sd136, 32'sd912,
32'sd1221, 32'sd175, 32'sd1624, 32'sd171, 32'sd1155, 32'sd1334,
32'sd1350, 32'sd179, 32'sd956, 32'sd1677, 32'sd1466, 32'sd753,
32'sd1665, 32'sd726, 32'sd684, 32'sd1448, 32'sd520, 32'sd679,
32'sd606, 32'sd1419, 32'sd1803, 32'sd836, 32'sd146, 32'sd1655,
32'sd828, 32'sd197, 32'sd1770, 32'sd313, 32'sd676, 32'sd139,
32'sd1516, 32'sd1409, 32'sd800, 32'sd1092, 32'sd1250, 32'sd1850,
32'sd1772, 32'sd683, 32'sd1053, 32'sd819, 32'sd1928, 32'sd1604,
32'sd1244, 32'sd975, 32'sd1192, 32'sd1180, 32'sd253, 32'sd1192,
32'sd272, 32'sd670, 32'sd1046, 32'sd1683, 32'sd1363, 32'sd1560,
32'sd1032, 32'sd1252, 32'sd524, 32'sd763, 32'sd739, 32'sd396,
32'sd171, 32'sd116, 32'sd1851, 32'sd217, 32'sd1247, 32'sd1858,
32'sd1092, 32'sd562, 32'sd544, 32'sd277, 32'sd593, 32'sd1673,
32'sd1457, 32'sd1603, 32'sd812, 32'sd1008, 32'sd1211, 32'sd1218,
32'sd1725, 32'sd556, 32'sd427, 32'sd1035, 32'sd647, 32'sd1943,
32'sd1229, 32'sd1123, 32'sd686, 32'sd1679, 32'sd754, 32'sd692,
32'sd594, 32'sd1115, 32'sd1507, 32'sd906, 32'sd1073, 32'sd1690,
32'sd1989, 32'sd1039, 32'sd935, 32'sd481, 32'sd1453, 32'sd1650,
32'sd463, 32'sd1209, 32'sd1330, 32'sd1549, 32'sd157, 32'sd1208,
32'sd1997, 32'sd1105, 32'sd304, 32'sd625, 32'sd1068, 32'sd1612,
32'sd1967, 32'sd874, 32'sd124, 32'sd1800, 32'sd685, 32'sd1360,
32'sd719, 32'sd1460, 32'sd1052, 32'sd1891, 32'sd207, 32'sd992,
32'sd1446, 32'sd949, 32'sd270, 32'sd716, 32'sd1650, 32'sd593,
32'sd362, 32'sd1611, 32'sd1830, 32'sd1724, 32'sd1042, 32'sd1023,
32'sd829, 32'sd1683, 32'sd1122, 32'sd862, 32'sd108, 32'sd280,
32'sd497, 32'sd654, 32'sd1445, 32'sd232, 32'sd1839, 32'sd1922,
32'sd1819, 32'sd1325, 32'sd1317, 32'sd657, 32'sd1409, 32'sd775,
32'sd826, 32'sd882, 32'sd1792, 32'sd710, 32'sd1850, 32'sd502,
32'sd630, 32'sd1011, 32'sd518, 32'sd1308, 32'sd851, 32'sd350,
32'sd941, 32'sd1788, 32'sd632, 32'sd790, 32'sd129, 32'sd1956,
32'sd928, 32'sd1837, 32'sd1745, 32'sd841, 32'sd1851, 32'sd1440,
32'sd1213, 32'sd1551, 32'sd278, 32'sd1833, 32'sd956, 32'sd666,
32'sd311, 32'sd739, 32'sd1034, 32'sd952, 32'sd1764, 32'sd1316,
32'sd1177, 32'sd1434, 32'sd1454, 32'sd603, 32'sd1092, 32'sd587,
32'sd408, 32'sd1532, 32'sd1846, 32'sd1605, 32'sd937, 32'sd971,
32'sd1507, 32'sd1703, 32'sd533, 32'sd463, 32'sd1165, 32'sd314,
32'sd1440, 32'sd1358, 32'sd1577, 32'sd1473, 32'sd1968, 32'sd341,
32'sd1983, 32'sd196, 32'sd934, 32'sd1980, 32'sd1631, 32'sd1574,
32'sd1157, 32'sd1365, 32'sd1859, 32'sd1975, 32'sd1036, 32'sd637,
32'sd1235, 32'sd1917, 32'sd1357, 32'sd1664, 32'sd283, 32'sd414,
32'sd967, 32'sd1006, 32'sd1319, 32'sd1606, 32'sd1867, 32'sd178,
32'sd144, 32'sd1464, 32'sd1311, 32'sd671, 32'sd328, 32'sd923,
32'sd785, 32'sd1950, 32'sd1393, 32'sd1584, 32'sd1440, 32'sd1576,
32'sd1713, 32'sd1878, 32'sd717, 32'sd743, 32'sd255, 32'sd227,
32'sd504, 32'sd1117, 32'sd1941, 32'sd1632, 32'sd626, 32'sd1430,
32'sd134, 32'sd406, 32'sd1376, 32'sd1522, 32'sd1780, 32'sd1217,
32'sd284, 32'sd1140, 32'sd1413, 32'sd1636, 32'sd755, 32'sd800,
32'sd180, 32'sd1775, 32'sd281, 32'sd1651, 32'sd419, 32'sd1224,
32'sd1879, 32'sd1861, 32'sd379, 32'sd325, 32'sd1637, 32'sd940,
32'sd1648, 32'sd1523, 32'sd306, 32'sd506, 32'sd380, 32'sd984,
32'sd953, 32'sd613, 32'sd1520, 32'sd967, 32'sd306, 32'sd836,
32'sd885, 32'sd378, 32'sd1530, 32'sd1873, 32'sd1604, 32'sd1279,
32'sd1151, 32'sd1637, 32'sd908, 32'sd1525, 32'sd1828, 32'sd1812,
32'sd1745, 32'sd966, 32'sd1418, 32'sd595, 32'sd1065, 32'sd1596,
32'sd595, 32'sd1435, 32'sd1109, 32'sd1842, 32'sd844, 32'sd1467,
32'sd1077, 32'sd944, 32'sd1338, 32'sd1024, 32'sd897, 32'sd1914,
32'sd1373, 32'sd559, 32'sd1951, 32'sd1424, 32'sd623, 32'sd1148,
32'sd103, 32'sd228, 32'sd1947, 32'sd1344, 32'sd1573, 32'sd1845,
32'sd685, 32'sd908, 32'sd1706, 32'sd707, 32'sd1552, 32'sd727,
32'sd435, 32'sd1120, 32'sd820, 32'sd325, 32'sd1168, 32'sd916,
32'sd205, 32'sd1054, 32'sd1644, 32'sd161, 32'sd948, 32'sd1686,
32'sd1424, 32'sd1228, 32'sd879, 32'sd566, 32'sd1211, 32'sd146,
32'sd1160, 32'sd465, 32'sd1944, 32'sd714, 32'sd1042, 32'sd803,
32'sd1969, 32'sd1345, 32'sd1135, 32'sd1866, 32'sd1819, 32'sd1516,
32'sd989, 32'sd376, 32'sd966, 32'sd440, 32'sd1924, 32'sd1549,
32'sd956, 32'sd607, 32'sd1277, 32'sd1460, 32'sd390, 32'sd1603,
32'sd120, 32'sd849, 32'sd989, 32'sd167, 32'sd1482, 32'sd1831,
32'sd1590, 32'sd650, 32'sd853, 32'sd185, 32'sd1954, 32'sd156,
32'sd949, 32'sd987, 32'sd406, 32'sd1252, 32'sd1464, 32'sd497,
32'sd136, 32'sd1629, 32'sd247, 32'sd1473, 32'sd915, 32'sd1919,
32'sd934, 32'sd942, 32'sd1949, 32'sd986, 32'sd1986, 32'sd678,
32'sd1352, 32'sd1561, 32'sd1342, 32'sd818, 32'sd1285, 32'sd1995,
32'sd1100, 32'sd1769, 32'sd1411, 32'sd1463, 32'sd938, 32'sd971,
32'sd1302, 32'sd473, 32'sd722, 32'sd1062, 32'sd875, 32'sd1460,
32'sd967, 32'sd584, 32'sd441, 32'sd406, 32'sd213, 32'sd433,
32'sd1361, 32'sd1281, 32'sd1153, 32'sd1423, 32'sd546, 32'sd958,
32'sd904, 32'sd781, 32'sd700, 32'sd1442, 32'sd294, 32'sd762,
32'sd1266, 32'sd1344, 32'sd170, 32'sd288, 32'sd1734, 32'sd823,
32'sd497, 32'sd149, 32'sd688, 32'sd542, 32'sd234, 32'sd490,
32'sd1397, 32'sd155, 32'sd1152, 32'sd807, 32'sd957, 32'sd462,
32'sd1765, 32'sd1265, 32'sd207, 32'sd1441, 32'sd1395, 32'sd1282,
32'sd343, 32'sd593, 32'sd410, 32'sd1727, 32'sd994, 32'sd1686,
32'sd530, 32'sd433, 32'sd1078, 32'sd1922, 32'sd400, 32'sd601,
32'sd303, 32'sd887, 32'sd471, 32'sd1809, 32'sd1690, 32'sd1516,
32'sd1125, 32'sd1028, 32'sd147, 32'sd862, 32'sd1184, 32'sd1604,
32'sd1557, 32'sd808, 32'sd1562, 32'sd1624, 32'sd1769, 32'sd567,
32'sd348, 32'sd437, 32'sd1233, 32'sd1665, 32'sd1200, 32'sd818,
32'sd1441, 32'sd435, 32'sd549, 32'sd1514, 32'sd792, 32'sd1328,
32'sd1916, 32'sd565, 32'sd1172, 32'sd1870, 32'sd1827, 32'sd1106,
32'sd1047, 32'sd690, 32'sd936, 32'sd1980, 32'sd954, 32'sd1204,
32'sd411, 32'sd696, 32'sd531, 32'sd1170, 32'sd1056, 32'sd341,
32'sd922, 32'sd1576, 32'sd1933, 32'sd1947, 32'sd1410, 32'sd278,
32'sd1849, 32'sd489, 32'sd1619, 32'sd621, 32'sd862, 32'sd1598,
32'sd1815, 32'sd1617, 32'sd1778, 32'sd1158, 32'sd518, 32'sd1134,
32'sd1551, 32'sd692, 32'sd1818, 32'sd1897, 32'sd409, 32'sd1765,
32'sd1894, 32'sd118, 32'sd1512, 32'sd172, 32'sd1092, 32'sd104,
32'sd1852, 32'sd103, 32'sd1291, 32'sd564, 32'sd1761, 32'sd1767,
32'sd158, 32'sd902, 32'sd1984, 32'sd562, 32'sd162, 32'sd1090,
32'sd1544, 32'sd1925, 32'sd563, 32'sd1382, 32'sd1511, 32'sd821,
32'sd326, 32'sd846, 32'sd889, 32'sd1447, 32'sd584, 32'sd1992,
32'sd202, 32'sd1911, 32'sd1566, 32'sd1889, 32'sd1115, 32'sd1887,
32'sd204, 32'sd429, 32'sd614, 32'sd1027, 32'sd1830, 32'sd1999,
32'sd978, 32'sd1132, 32'sd539, 32'sd660, 32'sd454, 32'sd939,
32'sd1193, 32'sd1479, 32'sd1866, 32'sd230, 32'sd1885, 32'sd628,
32'sd1937, 32'sd305, 32'sd1026, 32'sd129, 32'sd1108, 32'sd1852,
32'sd1984, 32'sd867, 32'sd1127, 32'sd411, 32'sd606, 32'sd624,
32'sd1533, 32'sd1588, 32'sd1188, 32'sd1281, 32'sd1833, 32'sd1674,
32'sd403, 32'sd726, 32'sd1981, 32'sd505, 32'sd1098, 32'sd289,
32'sd1514, 32'sd596, 32'sd1910, 32'sd683, 32'sd1797, 32'sd1668,
32'sd418, 32'sd670, 32'sd1740, 32'sd1779, 32'sd361, 32'sd1298,
32'sd319, 32'sd1118, 32'sd1699, 32'sd1969, 32'sd246, 32'sd167,
32'sd1121, 32'sd1222, 32'sd1164, 32'sd1584, 32'sd928, 32'sd310,
32'sd141, 32'sd846, 32'sd1091, 32'sd1474, 32'sd1979, 32'sd1860,
32'sd440, 32'sd1036, 32'sd604, 32'sd1468, 32'sd1184, 32'sd581,
32'sd1399, 32'sd1935, 32'sd1513, 32'sd302, 32'sd1293, 32'sd880,
32'sd230, 32'sd1507, 32'sd112, 32'sd492, 32'sd422, 32'sd1261,
32'sd1914, 32'sd1324, 32'sd1318, 32'sd611, 32'sd121, 32'sd1206,
32'sd759, 32'sd1383, 32'sd372, 32'sd1016, 32'sd490, 32'sd616,
32'sd1829, 32'sd239, 32'sd1459, 32'sd360, 32'sd1957, 32'sd1854,
32'sd1770, 32'sd1732, 32'sd714, 32'sd1639, 32'sd1602, 32'sd1483,
32'sd1486, 32'sd868, 32'sd1715, 32'sd856, 32'sd1775, 32'sd203,
32'sd1964, 32'sd1333, 32'sd1893, 32'sd288, 32'sd1715, 32'sd693,
32'sd804, 32'sd1087, 32'sd1170, 32'sd172, 32'sd1889, 32'sd481,
32'sd309, 32'sd1051, 32'sd1905, 32'sd1664, 32'sd1804, 32'sd1500,
32'sd1309, 32'sd1522, 32'sd1503, 32'sd490, 32'sd559, 32'sd448,
32'sd1927, 32'sd843, 32'sd1396, 32'sd1986, 32'sd1081, 32'sd1462,
32'sd633, 32'sd875, 32'sd592, 32'sd829, 32'sd1690, 32'sd1595,
32'sd610, 32'sd563, 32'sd1827, 32'sd389, 32'sd746, 32'sd870,
32'sd893, 32'sd1461, 32'sd1847, 32'sd429, 32'sd1484, 32'sd1051,
32'sd1712, 32'sd1332, 32'sd1852, 32'sd876, 32'sd1745, 32'sd1898,
32'sd1441, 32'sd886, 32'sd1168, 32'sd1945, 32'sd1236, 32'sd1509,
32'sd1229, 32'sd808, 32'sd1999, 32'sd556, 32'sd1986, 32'sd230,
32'sd1649, 32'sd621, 32'sd276, 32'sd482, 32'sd1010, 32'sd1869,
32'sd600, 32'sd888, 32'sd1338, 32'sd994, 32'sd1764, 32'sd1000,
32'sd1890, 32'sd1967, 32'sd553, 32'sd916, 32'sd1044, 32'sd534,
32'sd900, 32'sd1684, 32'sd1555, 32'sd493, 32'sd1998, 32'sd976,
32'sd126, 32'sd306, 32'sd943, 32'sd1248, 32'sd509, 32'sd211,
32'sd610, 32'sd1737, 32'sd1112, 32'sd1419, 32'sd701, 32'sd495,
32'sd414, 32'sd792, 32'sd980, 32'sd1727, 32'sd739, 32'sd259,
32'sd948, 32'sd1892, 32'sd1056, 32'sd1754, 32'sd1818, 32'sd475,
32'sd1568, 32'sd299, 32'sd1892, 32'sd195, 32'sd230, 32'sd1204,
32'sd1601, 32'sd391, 32'sd579, 32'sd1215, 32'sd1851, 32'sd414,
32'sd377, 32'sd1046, 32'sd1151, 32'sd492, 32'sd747, 32'sd1392,
32'sd1854, 32'sd633, 32'sd1042, 32'sd1127, 32'sd129, 32'sd1498,
32'sd1079, 32'sd1545, 32'sd1311, 32'sd504, 32'sd526, 32'sd1896,
32'sd1373, 32'sd1662, 32'sd251, 32'sd102, 32'sd1474, 32'sd271,
32'sd515, 32'sd107, 32'sd908, 32'sd997, 32'sd133, 32'sd361,
32'sd762, 32'sd1411, 32'sd336, 32'sd1238, 32'sd1105, 32'sd920,
32'sd441, 32'sd703, 32'sd690, 32'sd1360, 32'sd1030, 32'sd1124,
32'sd1718, 32'sd646, 32'sd1214, 32'sd816, 32'sd549, 32'sd1727,
32'sd656, 32'sd336, 32'sd630, 32'sd1453, 32'sd1360, 32'sd1375,
32'sd1079, 32'sd686, 32'sd1304, 32'sd1088, 32'sd658, 32'sd1355,
32'sd361, 32'sd1071, 32'sd306, 32'sd1457, 32'sd228, 32'sd703,
32'sd429, 32'sd1787, 32'sd963, 32'sd1928, 32'sd1541, 32'sd1049,
32'sd1759, 32'sd959, 32'sd786, 32'sd407, 32'sd146, 32'sd967,
32'sd651, 32'sd1536, 32'sd1249, 32'sd378, 32'sd1216, 32'sd108,
32'sd201, 32'sd1208, 32'sd238, 32'sd273, 32'sd1296, 32'sd1574,
32'sd295, 32'sd1985, 32'sd1022, 32'sd1808, 32'sd1274, 32'sd204,
32'sd706, 32'sd506, 32'sd1938, 32'sd374, 32'sd413, 32'sd1292,
32'sd1869, 32'sd711, 32'sd1213, 32'sd1104, 32'sd1091, 32'sd691,
32'sd1067, 32'sd136, 32'sd153, 32'sd1233, 32'sd1414, 32'sd348,
32'sd985, 32'sd121, 32'sd1194, 32'sd191, 32'sd484, 32'sd292,
32'sd434, 32'sd1659, 32'sd592, 32'sd994, 32'sd506, 32'sd1491,
32'sd1941, 32'sd783, 32'sd970, 32'sd1544, 32'sd751, 32'sd1444,
32'sd814, 32'sd658, 32'sd1341, 32'sd1219, 32'sd706, 32'sd243,
32'sd1897, 32'sd1785, 32'sd1262, 32'sd383, 32'sd327, 32'sd434,
32'sd701, 32'sd613, 32'sd1622, 32'sd1693, 32'sd1682, 32'sd155,
32'sd1025, 32'sd522, 32'sd110, 32'sd1758, 32'sd1454, 32'sd1429,
32'sd1950, 32'sd720, 32'sd341, 32'sd882, 32'sd1739, 32'sd1353,
32'sd1721, 32'sd752, 32'sd157, 32'sd575, 32'sd1272, 32'sd394,
32'sd1158, 32'sd204, 32'sd725, 32'sd1671, 32'sd529, 32'sd1905,
32'sd1234, 32'sd441, 32'sd203, 32'sd1348, 32'sd1549, 32'sd1282,
32'sd949, 32'sd150, 32'sd1687, 32'sd1603, 32'sd1025, 32'sd409,
32'sd657, 32'sd1124, 32'sd1688, 32'sd1883, 32'sd435, 32'sd1381,
32'sd1776, 32'sd524, 32'sd1294, 32'sd908, 32'sd1962, 32'sd614,
32'sd1289, 32'sd558, 32'sd828, 32'sd1971, 32'sd1122, 32'sd518,
32'sd1917, 32'sd151, 32'sd916, 32'sd394, 32'sd115, 32'sd1435,
32'sd1796, 32'sd754, 32'sd196, 32'sd1229, 32'sd883, 32'sd1292,
32'sd154, 32'sd401, 32'sd961, 32'sd986, 32'sd1406, 32'sd554,
32'sd141, 32'sd1799, 32'sd1563, 32'sd1516, 32'sd165, 32'sd1808,
32'sd1283, 32'sd1315, 32'sd1516, 32'sd1536, 32'sd1599, 32'sd1821,
32'sd301, 32'sd1816, 32'sd448, 32'sd717, 32'sd1780, 32'sd1152,
32'sd1853, 32'sd1619, 32'sd1821, 32'sd1139, 32'sd1483, 32'sd1359,
32'sd1955, 32'sd255, 32'sd871, 32'sd1612, 32'sd167, 32'sd1811,
32'sd1548, 32'sd595, 32'sd1758, 32'sd1317, 32'sd463, 32'sd251,
32'sd1106, 32'sd702, 32'sd355, 32'sd879, 32'sd1730, 32'sd1815,
32'sd627, 32'sd952, 32'sd1979, 32'sd1254, 32'sd541, 32'sd730,
32'sd1187, 32'sd1518, 32'sd1280, 32'sd1798, 32'sd684, 32'sd1720,
32'sd526, 32'sd274, 32'sd662, 32'sd1899, 32'sd361, 32'sd1447,
32'sd925, 32'sd1896, 32'sd1402, 32'sd1139, 32'sd1116, 32'sd1906,
32'sd838, 32'sd1775, 32'sd311, 32'sd1036, 32'sd1716, 32'sd1485,
32'sd1234, 32'sd793, 32'sd1498, 32'sd1666, 32'sd1188, 32'sd1163,
32'sd761, 32'sd1226, 32'sd1378, 32'sd1053, 32'sd257, 32'sd566,
32'sd1510, 32'sd790, 32'sd1873, 32'sd1843, 32'sd869, 32'sd193,
32'sd921, 32'sd1200, 32'sd279, 32'sd1319, 32'sd1033, 32'sd364,
32'sd1050, 32'sd357, 32'sd1682, 32'sd1643, 32'sd106, 32'sd1529,
32'sd1026, 32'sd1434, 32'sd964, 32'sd1608, 32'sd1026, 32'sd1816,
32'sd595, 32'sd1285, 32'sd186, 32'sd647, 32'sd252, 32'sd1972,
32'sd1183, 32'sd448, 32'sd720, 32'sd883, 32'sd1801, 32'sd918,
32'sd786, 32'sd509, 32'sd545, 32'sd1521, 32'sd431, 32'sd1181,
32'sd1840, 32'sd686, 32'sd455, 32'sd796, 32'sd1680, 32'sd1684,
32'sd1463, 32'sd1163, 32'sd1010, 32'sd348, 32'sd870, 32'sd1648,
32'sd1518, 32'sd1750, 32'sd915, 32'sd1759, 32'sd1593, 32'sd651,
32'sd1081, 32'sd214, 32'sd320, 32'sd700, 32'sd1524, 32'sd285,
32'sd734, 32'sd1082, 32'sd887, 32'sd1063, 32'sd627, 32'sd1982,
32'sd1995, 32'sd199, 32'sd350, 32'sd508, 32'sd1598, 32'sd1959,
32'sd1653, 32'sd1038, 32'sd1057, 32'sd657, 32'sd1542, 32'sd1527,
32'sd1067, 32'sd1917, 32'sd1453, 32'sd259, 32'sd839, 32'sd246,
32'sd1837, 32'sd1944, 32'sd986, 32'sd1257, 32'sd1185, 32'sd1829,
32'sd560, 32'sd1519, 32'sd824, 32'sd627, 32'sd1491, 32'sd889,
32'sd1166, 32'sd1236, 32'sd1267, 32'sd583, 32'sd1746, 32'sd319,
32'sd1088, 32'sd1390, 32'sd1312, 32'sd1879, 32'sd958, 32'sd1662,
32'sd1118, 32'sd767, 32'sd387, 32'sd1669, 32'sd182, 32'sd1753,
32'sd783, 32'sd1930, 32'sd1335, 32'sd599, 32'sd1215, 32'sd1164,
32'sd1216, 32'sd1633, 32'sd278, 32'sd1243, 32'sd1348, 32'sd1389,
32'sd1951, 32'sd705, 32'sd1284, 32'sd1210, 32'sd1862, 32'sd773,
32'sd1466, 32'sd1234, 32'sd443, 32'sd1427, 32'sd122, 32'sd719,
32'sd1090, 32'sd202, 32'sd993, 32'sd1618, 32'sd257, 32'sd913,
32'sd1161, 32'sd283, 32'sd376, 32'sd963, 32'sd1478, 32'sd795,
32'sd1847, 32'sd1613, 32'sd343, 32'sd1021, 32'sd1765, 32'sd624,
32'sd897, 32'sd1868, 32'sd569, 32'sd660, 32'sd1243, 32'sd486,
32'sd238, 32'sd927, 32'sd1408, 32'sd1145, 32'sd184, 32'sd1808,
32'sd589, 32'sd1663, 32'sd278, 32'sd1826, 32'sd774, 32'sd1442,
32'sd1627, 32'sd1398, 32'sd885, 32'sd1611, 32'sd1326, 32'sd1189,
32'sd1913, 32'sd1343, 32'sd135, 32'sd281, 32'sd319, 32'sd535,
32'sd458, 32'sd1065, 32'sd783, 32'sd1273, 32'sd1913, 32'sd483,
32'sd446, 32'sd1207, 32'sd1930, 32'sd1911, 32'sd1501, 32'sd246,
32'sd1665, 32'sd112, 32'sd1831, 32'sd1659, 32'sd838, 32'sd252,
32'sd1472, 32'sd289, 32'sd1402, 32'sd1747, 32'sd753, 32'sd641,
32'sd408, 32'sd685, 32'sd138, 32'sd1605, 32'sd1307, 32'sd1649,
32'sd1488, 32'sd1659, 32'sd406, 32'sd350, 32'sd1372, 32'sd651,
32'sd1700, 32'sd1940, 32'sd1905, 32'sd530, 32'sd868, 32'sd175,
32'sd170, 32'sd1765, 32'sd1783, 32'sd1932, 32'sd720, 32'sd360,
32'sd1817, 32'sd430, 32'sd1920, 32'sd1669, 32'sd356, 32'sd784,
32'sd1131, 32'sd988, 32'sd1459, 32'sd1786, 32'sd1197, 32'sd645,
32'sd656, 32'sd800, 32'sd761, 32'sd1740, 32'sd1756, 32'sd757,
32'sd827, 32'sd264, 32'sd137, 32'sd1905, 32'sd1507, 32'sd1676,
32'sd1244, 32'sd1387, 32'sd251, 32'sd566, 32'sd1293, 32'sd119,
32'sd1157, 32'sd1393, 32'sd1386, 32'sd1334, 32'sd575, 32'sd1228,
32'sd866, 32'sd314, 32'sd1996, 32'sd1204, 32'sd1894, 32'sd1936,
32'sd860, 32'sd1036, 32'sd611, 32'sd732, 32'sd422, 32'sd846,
32'sd1133, 32'sd236, 32'sd1468, 32'sd828, 32'sd536, 32'sd306,
32'sd954, 32'sd823, 32'sd1166, 32'sd341, 32'sd1715, 32'sd266,
32'sd563, 32'sd1208, 32'sd1966, 32'sd1070, 32'sd1799, 32'sd1398,
32'sd1782, 32'sd595, 32'sd1406, 32'sd103, 32'sd391, 32'sd1245,
32'sd747, 32'sd1361, 32'sd1084, 32'sd1560, 32'sd1741, 32'sd1471,
32'sd270, 32'sd839, 32'sd1989, 32'sd911, 32'sd757, 32'sd672,
32'sd846, 32'sd1497, 32'sd216, 32'sd165, 32'sd295, 32'sd438,
32'sd1832, 32'sd1220, 32'sd1555, 32'sd1698, 32'sd186, 32'sd460,
32'sd312, 32'sd1352, 32'sd731, 32'sd1978, 32'sd1416, 32'sd1046,
32'sd165, 32'sd1152, 32'sd1087, 32'sd541, 32'sd1844, 32'sd1072,
32'sd510, 32'sd667, 32'sd121, 32'sd1377, 32'sd1242, 32'sd1013,
32'sd1384, 32'sd1421, 32'sd868, 32'sd295, 32'sd216, 32'sd747,
32'sd1452, 32'sd653, 32'sd1190, 32'sd1363, 32'sd636, 32'sd883,
32'sd716, 32'sd640, 32'sd1977, 32'sd1140, 32'sd1887, 32'sd1614,
32'sd737, 32'sd1268, 32'sd938, 32'sd960, 32'sd1677, 32'sd924,
32'sd327, 32'sd156, 32'sd1058, 32'sd386, 32'sd496, 32'sd286,
32'sd613, 32'sd683, 32'sd1155, 32'sd845, 32'sd132, 32'sd1573,
32'sd1607, 32'sd1776, 32'sd365, 32'sd1557, 32'sd1234, 32'sd884,
32'sd271, 32'sd1740, 32'sd586, 32'sd2000, 32'sd1010, 32'sd345,
32'sd784, 32'sd547, 32'sd1487, 32'sd401, 32'sd689, 32'sd1645,
32'sd1338, 32'sd349, 32'sd1809, 32'sd1306, 32'sd798, 32'sd1115,
32'sd1422, 32'sd820, 32'sd1893, 32'sd464, 32'sd376, 32'sd1713,
32'sd1996, 32'sd1660, 32'sd1455, 32'sd925, 32'sd1356, 32'sd836,
32'sd933, 32'sd1607, 32'sd1586, 32'sd1934, 32'sd745, 32'sd1757,
32'sd1713, 32'sd1634, 32'sd1230, 32'sd1863, 32'sd1906, 32'sd419,
32'sd1128, 32'sd1189, 32'sd1346, 32'sd1127, 32'sd678, 32'sd1759,
32'sd398, 32'sd645, 32'sd802, 32'sd1908, 32'sd1057, 32'sd1664,
32'sd657, 32'sd1254, 32'sd1071, 32'sd1825, 32'sd809, 32'sd1685,
32'sd1996, 32'sd1061, 32'sd993, 32'sd1240, 32'sd900, 32'sd385,
32'sd878, 32'sd1878, 32'sd1905, 32'sd1246, 32'sd1638, 32'sd116,
32'sd1857, 32'sd1417, 32'sd1054, 32'sd1714, 32'sd1872, 32'sd1276,
32'sd557, 32'sd1428, 32'sd1035, 32'sd1866, 32'sd118, 32'sd766,
32'sd1160, 32'sd1478, 32'sd1954, 32'sd472, 32'sd1676, 32'sd1106,
32'sd935, 32'sd1099, 32'sd1239, 32'sd378, 32'sd1674, 32'sd924,
32'sd1781, 32'sd306, 32'sd964, 32'sd1789, 32'sd1891, 32'sd1203,
32'sd1167, 32'sd352, 32'sd1939, 32'sd121, 32'sd1668, 32'sd1122,
32'sd1269, 32'sd1127, 32'sd273, 32'sd173, 32'sd172, 32'sd1793,
32'sd1110, 32'sd486, 32'sd1581, 32'sd1586, 32'sd1804, 32'sd742,
32'sd1220, 32'sd1958, 32'sd681, 32'sd1474, 32'sd976, 32'sd1540,
32'sd492, 32'sd694, 32'sd1821, 32'sd1254, 32'sd409, 32'sd321,
32'sd1719, 32'sd1127, 32'sd1657, 32'sd1395, 32'sd843, 32'sd1626,
32'sd104, 32'sd247, 32'sd1273, 32'sd1041, 32'sd731, 32'sd127,
32'sd864, 32'sd1919, 32'sd129, 32'sd444, 32'sd1357, 32'sd1184,
32'sd1356, 32'sd256, 32'sd1001, 32'sd1291, 32'sd647, 32'sd802,
32'sd1386, 32'sd1833, 32'sd182, 32'sd773, 32'sd1500, 32'sd1249,
32'sd243, 32'sd1084, 32'sd1151, 32'sd432, 32'sd124, 32'sd499,
32'sd1967, 32'sd1339, 32'sd1793, 32'sd1829, 32'sd713, 32'sd1553,
32'sd775, 32'sd183, 32'sd1922, 32'sd917, 32'sd288, 32'sd374,
32'sd1307, 32'sd1647, 32'sd1958, 32'sd596, 32'sd480, 32'sd1850,
32'sd1065, 32'sd1124, 32'sd1713, 32'sd1731, 32'sd1530, 32'sd1191,
32'sd1929, 32'sd413, 32'sd622, 32'sd1049, 32'sd1578, 32'sd1699,
32'sd1478, 32'sd1842, 32'sd1316, 32'sd1516, 32'sd830, 32'sd1079,
32'sd1867, 32'sd114, 32'sd1575, 32'sd1780, 32'sd160, 32'sd1124,
32'sd321, 32'sd879, 32'sd1161, 32'sd1579, 32'sd1332, 32'sd1071,
32'sd385, 32'sd1652, 32'sd793, 32'sd1539, 32'sd1301, 32'sd214,
32'sd1551, 32'sd1419, 32'sd1861, 32'sd666, 32'sd1720, 32'sd295,
32'sd1841, 32'sd1420, 32'sd866, 32'sd475, 32'sd1312, 32'sd872,
32'sd518, 32'sd1156, 32'sd680, 32'sd185, 32'sd1718, 32'sd756,
32'sd1315, 32'sd1272, 32'sd1950, 32'sd1578, 32'sd196, 32'sd1733,
32'sd1618, 32'sd1863, 32'sd707, 32'sd824, 32'sd1397, 32'sd1889,
32'sd1563, 32'sd1787, 32'sd984, 32'sd1937, 32'sd1646, 32'sd1004,
32'sd728, 32'sd1994, 32'sd1719, 32'sd1236, 32'sd1878, 32'sd1148,
32'sd175, 32'sd558, 32'sd1699, 32'sd181, 32'sd1168, 32'sd937,
32'sd321, 32'sd1987, 32'sd577, 32'sd1825, 32'sd219, 32'sd128,
32'sd426, 32'sd615, 32'sd639, 32'sd713, 32'sd701, 32'sd1935,
32'sd605, 32'sd1106, 32'sd1265, 32'sd167, 32'sd321, 32'sd1562,
32'sd1705, 32'sd209, 32'sd285, 32'sd985, 32'sd1631, 32'sd444,
32'sd1670, 32'sd141, 32'sd711, 32'sd466, 32'sd1181, 32'sd755,
32'sd565, 32'sd427, 32'sd376, 32'sd1515, 32'sd1403, 32'sd1847,
32'sd191, 32'sd1231, 32'sd137, 32'sd1341, 32'sd1700, 32'sd1236,
32'sd225, 32'sd306, 32'sd1282, 32'sd1069, 32'sd419, 32'sd417,
32'sd972, 32'sd1719, 32'sd1770, 32'sd1689, 32'sd968, 32'sd1418,
32'sd269, 32'sd1755, 32'sd689, 32'sd372, 32'sd883, 32'sd1793,
32'sd1840, 32'sd1999, 32'sd433, 32'sd1361, 32'sd1066, 32'sd292,
32'sd376, 32'sd1049, 32'sd1847, 32'sd146, 32'sd1686, 32'sd920,
32'sd1441, 32'sd1621, 32'sd1380, 32'sd146, 32'sd1208, 32'sd927,
32'sd1775, 32'sd324, 32'sd494, 32'sd298, 32'sd902, 32'sd1495,
32'sd887, 32'sd1927, 32'sd121, 32'sd774, 32'sd429, 32'sd349,
32'sd1595, 32'sd1374, 32'sd1871, 32'sd271, 32'sd359, 32'sd510,
32'sd1713, 32'sd918, 32'sd862, 32'sd758, 32'sd1637, 32'sd1429,
32'sd1565, 32'sd1437, 32'sd984, 32'sd131, 32'sd236, 32'sd305,
32'sd1139, 32'sd746, 32'sd1342, 32'sd1554, 32'sd1549, 32'sd1550,
32'sd1624, 32'sd596, 32'sd546, 32'sd999, 32'sd1913, 32'sd1651,
32'sd1312, 32'sd888, 32'sd580, 32'sd1259, 32'sd1237, 32'sd1508,
32'sd171, 32'sd265, 32'sd1006, 32'sd788, 32'sd222, 32'sd472,
32'sd357, 32'sd1770, 32'sd1590, 32'sd1809, 32'sd1243, 32'sd1034,
32'sd443, 32'sd907, 32'sd335, 32'sd1832, 32'sd412, 32'sd1087,
32'sd1862, 32'sd1947, 32'sd1586, 32'sd315, 32'sd1758, 32'sd142,
32'sd1609, 32'sd1774, 32'sd1751, 32'sd531, 32'sd320, 32'sd1606,
32'sd1064, 32'sd1402, 32'sd1663, 32'sd1789, 32'sd1471, 32'sd323,
32'sd838, 32'sd1615, 32'sd548, 32'sd633, 32'sd1388, 32'sd799,
32'sd1539, 32'sd1427, 32'sd336, 32'sd1607, 32'sd329, 32'sd1695,
32'sd697, 32'sd207, 32'sd1459, 32'sd288, 32'sd1607, 32'sd1157,
32'sd580, 32'sd1874, 32'sd286, 32'sd1967, 32'sd1613, 32'sd1965,
32'sd544, 32'sd997, 32'sd1507, 32'sd106, 32'sd1766, 32'sd536,
32'sd1860, 32'sd1014, 32'sd1216, 32'sd1992, 32'sd385, 32'sd1665,
32'sd515, 32'sd1157, 32'sd1836, 32'sd1638, 32'sd1072, 32'sd1331,
32'sd508, 32'sd191, 32'sd130, 32'sd1151, 32'sd514, 32'sd589,
32'sd1642, 32'sd463, 32'sd172, 32'sd189, 32'sd587, 32'sd1598,
32'sd1231, 32'sd1225, 32'sd1184, 32'sd838, 32'sd1046, 32'sd1147,
32'sd1650, 32'sd1550, 32'sd1212, 32'sd1378, 32'sd778, 32'sd1737,
32'sd1760, 32'sd1526, 32'sd1416, 32'sd1594, 32'sd1078, 32'sd1746,
32'sd302, 32'sd1357, 32'sd1626, 32'sd1123, 32'sd1090, 32'sd416,
32'sd1670, 32'sd168, 32'sd854, 32'sd702, 32'sd993, 32'sd535,
32'sd1900, 32'sd659, 32'sd678, 32'sd1663, 32'sd1246, 32'sd1371,
32'sd973, 32'sd488, 32'sd276, 32'sd800, 32'sd833, 32'sd1411,
32'sd1477, 32'sd1953, 32'sd1689, 32'sd1596, 32'sd1965, 32'sd701,
32'sd1395, 32'sd177, 32'sd218, 32'sd295, 32'sd1504, 32'sd124,
32'sd776, 32'sd383, 32'sd1117, 32'sd517, 32'sd872, 32'sd915,
32'sd259, 32'sd1856, 32'sd1060, 32'sd491, 32'sd132, 32'sd336,
32'sd1882, 32'sd480, 32'sd587, 32'sd1101, 32'sd229, 32'sd1496,
32'sd1853, 32'sd1144, 32'sd325, 32'sd1275, 32'sd979, 32'sd840,
32'sd1066, 32'sd1465, 32'sd1330, 32'sd571, 32'sd189, 32'sd345,
32'sd115, 32'sd138, 32'sd133, 32'sd1355, 32'sd1580, 32'sd1698,
32'sd1726, 32'sd1562, 32'sd320, 32'sd231, 32'sd1605, 32'sd916,
32'sd1558, 32'sd644, 32'sd1341, 32'sd1933, 32'sd1918, 32'sd760,
32'sd752, 32'sd912, 32'sd592, 32'sd1939, 32'sd529, 32'sd642,
32'sd1947, 32'sd923, 32'sd382, 32'sd1243, 32'sd1493, 32'sd184,
32'sd1772, 32'sd1989, 32'sd676, 32'sd1655, 32'sd1163, 32'sd561,
32'sd806, 32'sd735, 32'sd1985, 32'sd1273, 32'sd1681, 32'sd1471,
32'sd1200, 32'sd1609, 32'sd408, 32'sd766, 32'sd1498, 32'sd786,
32'sd562, 32'sd1001, 32'sd1565, 32'sd1275, 32'sd785, 32'sd589,
32'sd677, 32'sd317, 32'sd1987, 32'sd663, 32'sd156, 32'sd1166,
32'sd960, 32'sd1189, 32'sd145, 32'sd379, 32'sd863, 32'sd1807,
32'sd1912, 32'sd382, 32'sd1299, 32'sd203, 32'sd1488, 32'sd1006,
32'sd641, 32'sd594, 32'sd921, 32'sd1096, 32'sd1231, 32'sd1244,
32'sd398, 32'sd1649, 32'sd159, 32'sd1375, 32'sd907, 32'sd601,
32'sd346, 32'sd302, 32'sd797, 32'sd1208, 32'sd104, 32'sd522,
32'sd1212, 32'sd432, 32'sd920, 32'sd198, 32'sd1235, 32'sd1742,
32'sd412, 32'sd1792, 32'sd1773, 32'sd1590, 32'sd143, 32'sd310,
32'sd284, 32'sd1377, 32'sd588, 32'sd809, 32'sd794, 32'sd535,
32'sd312, 32'sd530, 32'sd313, 32'sd126, 32'sd676, 32'sd1483,
32'sd487, 32'sd177, 32'sd264, 32'sd1953, 32'sd802, 32'sd1943,
32'sd1549, 32'sd1126, 32'sd308, 32'sd1004, 32'sd711, 32'sd1677,
32'sd1758, 32'sd774, 32'sd1685, 32'sd913, 32'sd1917, 32'sd1529,
32'sd1216, 32'sd1138, 32'sd1685, 32'sd1707, 32'sd550, 32'sd1546,
32'sd1359, 32'sd457, 32'sd441, 32'sd1129, 32'sd239, 32'sd824,
32'sd725, 32'sd897, 32'sd1440, 32'sd524, 32'sd599, 32'sd978,
32'sd487, 32'sd1960, 32'sd217, 32'sd646, 32'sd838, 32'sd1222,
32'sd1175, 32'sd1083, 32'sd1686, 32'sd365, 32'sd1730, 32'sd684,
32'sd159, 32'sd104, 32'sd359, 32'sd1366, 32'sd1899, 32'sd176,
32'sd1186, 32'sd1295, 32'sd1353, 32'sd1625, 32'sd1540, 32'sd1867,
32'sd920, 32'sd1131, 32'sd164, 32'sd164, 32'sd1788, 32'sd1379,
32'sd1844, 32'sd618, 32'sd928, 32'sd1738, 32'sd1344, 32'sd526,
32'sd538, 32'sd1219, 32'sd230, 32'sd567, 32'sd1074, 32'sd458,
32'sd1760, 32'sd1179, 32'sd397, 32'sd849, 32'sd119, 32'sd1924,
32'sd1741, 32'sd335, 32'sd738, 32'sd318, 32'sd493, 32'sd1739,
32'sd129, 32'sd764, 32'sd616, 32'sd689, 32'sd557, 32'sd1965,
32'sd1828, 32'sd154, 32'sd1250, 32'sd434, 32'sd535, 32'sd490,
32'sd1549, 32'sd1315, 32'sd138, 32'sd960, 32'sd1049, 32'sd1554,
32'sd1000, 32'sd1637, 32'sd378, 32'sd1057, 32'sd1751, 32'sd1401,
32'sd407, 32'sd1002, 32'sd1668, 32'sd383, 32'sd1390, 32'sd1634,
32'sd1201, 32'sd1646, 32'sd1046, 32'sd612, 32'sd572, 32'sd613,
32'sd135, 32'sd1747, 32'sd364, 32'sd822, 32'sd1416, 32'sd1887,
32'sd1236, 32'sd1886, 32'sd1351, 32'sd507, 32'sd1971, 32'sd1479,
32'sd1819, 32'sd1690, 32'sd1481, 32'sd409, 32'sd439, 32'sd860,
32'sd350, 32'sd223, 32'sd1642, 32'sd199, 32'sd1413, 32'sd1916,
32'sd624, 32'sd270, 32'sd1917, 32'sd1008, 32'sd832, 32'sd384,
32'sd1008, 32'sd248, 32'sd1483, 32'sd121, 32'sd1749, 32'sd1087,
32'sd1735, 32'sd1432, 32'sd200, 32'sd1141, 32'sd1609, 32'sd1812,
32'sd1397, 32'sd1369, 32'sd223, 32'sd903, 32'sd1692, 32'sd822,
32'sd251, 32'sd1739, 32'sd1268, 32'sd1329, 32'sd157, 32'sd284,
32'sd1183, 32'sd1950, 32'sd933, 32'sd976, 32'sd1280, 32'sd1236,
32'sd1404, 32'sd452, 32'sd750, 32'sd1319, 32'sd125, 32'sd1097,
32'sd701, 32'sd1099, 32'sd500, 32'sd897, 32'sd1145, 32'sd1173,
32'sd1292, 32'sd438, 32'sd1756, 32'sd1429, 32'sd971, 32'sd356,
32'sd1401, 32'sd267, 32'sd1491, 32'sd1923, 32'sd972, 32'sd1283,
32'sd642, 32'sd1499, 32'sd1775, 32'sd1951, 32'sd1504, 32'sd816,
32'sd666, 32'sd1462, 32'sd656, 32'sd134, 32'sd351, 32'sd468,
32'sd918, 32'sd736, 32'sd132, 32'sd1003, 32'sd1022, 32'sd1516,
32'sd1917, 32'sd1288, 32'sd122, 32'sd1769, 32'sd1276, 32'sd831,
32'sd554, 32'sd218, 32'sd932, 32'sd1707, 32'sd451, 32'sd1082,
32'sd1474, 32'sd447, 32'sd1863, 32'sd315, 32'sd1733, 32'sd1245,
32'sd853, 32'sd517, 32'sd1763, 32'sd1552, 32'sd307, 32'sd966,
32'sd637, 32'sd1744, 32'sd608, 32'sd804, 32'sd1220, 32'sd273,
32'sd540, 32'sd1134, 32'sd1744, 32'sd114, 32'sd1938, 32'sd961,
32'sd313, 32'sd793, 32'sd989, 32'sd1470, 32'sd284, 32'sd1829,
32'sd1622, 32'sd1648, 32'sd394, 32'sd236, 32'sd764, 32'sd682,
32'sd341, 32'sd820, 32'sd699, 32'sd136, 32'sd328, 32'sd1360,
32'sd1807, 32'sd1275, 32'sd1802, 32'sd1360, 32'sd814, 32'sd672,
32'sd1723, 32'sd1361, 32'sd954, 32'sd361, 32'sd1285, 32'sd526,
32'sd1101, 32'sd124, 32'sd445, 32'sd1528, 32'sd1115, 32'sd546,
32'sd548, 32'sd1173, 32'sd1554, 32'sd645, 32'sd308, 32'sd1425,
32'sd1552, 32'sd1312, 32'sd784, 32'sd1628, 32'sd406, 32'sd1015,
32'sd829, 32'sd204, 32'sd352, 32'sd1785, 32'sd216, 32'sd1031,
32'sd1276, 32'sd815, 32'sd1046, 32'sd1676, 32'sd1713, 32'sd145,
32'sd1459, 32'sd434, 32'sd767, 32'sd711, 32'sd1389, 32'sd368,
32'sd1808, 32'sd610, 32'sd331, 32'sd720, 32'sd160, 32'sd1854,
32'sd912, 32'sd1455, 32'sd435, 32'sd916, 32'sd1324, 32'sd222,
32'sd450, 32'sd1270, 32'sd860, 32'sd1752, 32'sd1200, 32'sd645,
32'sd1866, 32'sd1324, 32'sd1551, 32'sd999, 32'sd659, 32'sd580,
32'sd1716, 32'sd1782, 32'sd1225, 32'sd997, 32'sd658, 32'sd1197,
32'sd217, 32'sd786, 32'sd657, 32'sd1567, 32'sd1652, 32'sd238,
32'sd1940, 32'sd267, 32'sd196, 32'sd768, 32'sd1176, 32'sd1526,
32'sd1721, 32'sd804, 32'sd474, 32'sd312, 32'sd1066, 32'sd196,
32'sd781, 32'sd809, 32'sd373, 32'sd816, 32'sd1915, 32'sd679,
32'sd1139, 32'sd943, 32'sd1987, 32'sd1128, 32'sd822, 32'sd1214,
32'sd306, 32'sd924, 32'sd635, 32'sd444, 32'sd273, 32'sd181,
32'sd926, 32'sd1968, 32'sd1222, 32'sd860, 32'sd1406, 32'sd1292,
32'sd906, 32'sd1298, 32'sd220, 32'sd1519, 32'sd792, 32'sd1765,
32'sd1304, 32'sd1505, 32'sd1549, 32'sd271, 32'sd103, 32'sd386,
32'sd1832, 32'sd1649, 32'sd1737, 32'sd720, 32'sd567, 32'sd1549,
32'sd1914, 32'sd1917, 32'sd993, 32'sd1426, 32'sd1497, 32'sd1101,
32'sd1250, 32'sd1864, 32'sd179, 32'sd1742, 32'sd1027, 32'sd434,
32'sd1949, 32'sd1996, 32'sd1290, 32'sd1563, 32'sd1186, 32'sd1456,
32'sd1823, 32'sd1828, 32'sd1034, 32'sd935, 32'sd1759, 32'sd712,
32'sd283, 32'sd351, 32'sd1586, 32'sd853, 32'sd481, 32'sd1084,
32'sd1933, 32'sd1312, 32'sd934, 32'sd319, 32'sd1224, 32'sd1204,
32'sd1126, 32'sd1365, 32'sd887, 32'sd1782, 32'sd1592, 32'sd1199,
32'sd122, 32'sd1871, 32'sd1462, 32'sd1616, 32'sd417, 32'sd1267,
32'sd1035, 32'sd844, 32'sd1720, 32'sd1605, 32'sd365, 32'sd1910,
32'sd1284, 32'sd200, 32'sd909, 32'sd348, 32'sd528, 32'sd1861,
32'sd207, 32'sd466, 32'sd1513, 32'sd531, 32'sd817, 32'sd423,
32'sd1139, 32'sd1982, 32'sd1329, 32'sd1496, 32'sd444, 32'sd1909,
32'sd553, 32'sd214, 32'sd375, 32'sd320, 32'sd406, 32'sd1201,
32'sd259, 32'sd1805, 32'sd808, 32'sd226, 32'sd223, 32'sd1724,
32'sd414, 32'sd910, 32'sd1399, 32'sd781, 32'sd1945, 32'sd143,
32'sd1528, 32'sd1991, 32'sd990, 32'sd1443, 32'sd1098, 32'sd1769,
32'sd1908, 32'sd1359, 32'sd320, 32'sd1782, 32'sd473, 32'sd1944,
32'sd1319, 32'sd598, 32'sd146, 32'sd1758, 32'sd222, 32'sd1183,
32'sd1600, 32'sd374, 32'sd1994, 32'sd724, 32'sd658, 32'sd1931,
32'sd697, 32'sd117, 32'sd305, 32'sd883, 32'sd1681, 32'sd1844,
32'sd632, 32'sd827, 32'sd1386, 32'sd1454, 32'sd486, 32'sd1165,
32'sd1891, 32'sd1177, 32'sd691, 32'sd853, 32'sd1329, 32'sd1058,
32'sd1517, 32'sd1319, 32'sd343, 32'sd1040, 32'sd1691, 32'sd790,
32'sd1039, 32'sd1068, 32'sd782, 32'sd1510, 32'sd219, 32'sd291,
32'sd1257, 32'sd492, 32'sd1845, 32'sd1328, 32'sd719, 32'sd431,
32'sd713, 32'sd907, 32'sd1155, 32'sd1839, 32'sd1125, 32'sd1908,
32'sd1760, 32'sd256, 32'sd1024, 32'sd1496, 32'sd1762, 32'sd1150,
32'sd837, 32'sd588, 32'sd466, 32'sd512, 32'sd699, 32'sd1758,
32'sd1963, 32'sd1548, 32'sd388, 32'sd1591, 32'sd462, 32'sd757,
32'sd1457, 32'sd507, 32'sd696, 32'sd734, 32'sd392, 32'sd1713,
32'sd1042, 32'sd1529, 32'sd1948, 32'sd449, 32'sd1138, 32'sd543,
32'sd706, 32'sd479, 32'sd699, 32'sd1332, 32'sd1802, 32'sd1297,
32'sd968, 32'sd909, 32'sd320, 32'sd625, 32'sd240, 32'sd140,
32'sd1076, 32'sd105, 32'sd1548, 32'sd1616, 32'sd167, 32'sd195,
32'sd933, 32'sd1817, 32'sd1401, 32'sd1160, 32'sd299, 32'sd297,
32'sd154, 32'sd601, 32'sd1645, 32'sd1419, 32'sd597, 32'sd1623,
32'sd1956, 32'sd700, 32'sd1979, 32'sd1786, 32'sd116, 32'sd1450,
32'sd958, 32'sd1297, 32'sd1890, 32'sd1895, 32'sd576, 32'sd990,
32'sd1929, 32'sd1292, 32'sd203, 32'sd1523, 32'sd187, 32'sd585,
32'sd1965, 32'sd1041, 32'sd1517, 32'sd673, 32'sd436, 32'sd605,
32'sd1417, 32'sd366, 32'sd1745, 32'sd1525, 32'sd1902, 32'sd1866,
32'sd1965, 32'sd122, 32'sd495, 32'sd561, 32'sd143, 32'sd1818,
32'sd1987, 32'sd1461, 32'sd1375, 32'sd1099, 32'sd1089, 32'sd1701,
32'sd1512, 32'sd500, 32'sd800, 32'sd1072, 32'sd1581, 32'sd469,
32'sd182, 32'sd1299, 32'sd617, 32'sd195, 32'sd1876, 32'sd1589,
32'sd119, 32'sd1159, 32'sd350, 32'sd1993, 32'sd1492, 32'sd212,
32'sd1966, 32'sd602, 32'sd622, 32'sd1495, 32'sd1584, 32'sd786,
32'sd1762, 32'sd744, 32'sd798, 32'sd525, 32'sd112, 32'sd1390,
32'sd1405, 32'sd1384, 32'sd1680, 32'sd1123, 32'sd172, 32'sd570,
32'sd1662, 32'sd455, 32'sd1867, 32'sd697, 32'sd749, 32'sd1622,
32'sd940, 32'sd1640, 32'sd1988, 32'sd1393, 32'sd595, 32'sd1482,
32'sd1351, 32'sd1570, 32'sd1905, 32'sd467, 32'sd374, 32'sd432,
32'sd459, 32'sd691, 32'sd1469, 32'sd1492, 32'sd879, 32'sd1692,
32'sd1896, 32'sd1113, 32'sd1233, 32'sd1867, 32'sd1405, 32'sd1055,
32'sd259, 32'sd1533, 32'sd1936, 32'sd685, 32'sd1846, 32'sd266,
32'sd1388, 32'sd937, 32'sd1257, 32'sd1709, 32'sd1330, 32'sd1792,
32'sd558, 32'sd612, 32'sd1380, 32'sd876, 32'sd191, 32'sd1689,
32'sd1662, 32'sd437, 32'sd588, 32'sd206, 32'sd1813, 32'sd1753,
32'sd380, 32'sd1218, 32'sd754, 32'sd617, 32'sd1247, 32'sd1079,
32'sd239, 32'sd406, 32'sd520, 32'sd349, 32'sd753, 32'sd1147,
32'sd209, 32'sd1559, 32'sd801, 32'sd419, 32'sd1958, 32'sd1091,
32'sd664, 32'sd1526, 32'sd183, 32'sd1310, 32'sd1793, 32'sd1559,
32'sd975, 32'sd888, 32'sd972, 32'sd354, 32'sd972, 32'sd575,
32'sd420, 32'sd1846, 32'sd1592, 32'sd1334, 32'sd307, 32'sd1992,
32'sd591, 32'sd877, 32'sd904, 32'sd334, 32'sd967, 32'sd1835,
32'sd1106, 32'sd1871, 32'sd288, 32'sd1651, 32'sd1107, 32'sd1498,
32'sd1097, 32'sd1242, 32'sd420, 32'sd1534, 32'sd622, 32'sd669,
32'sd346, 32'sd1073, 32'sd1006, 32'sd1418, 32'sd704, 32'sd1433,
32'sd1883, 32'sd1467, 32'sd1738, 32'sd1822, 32'sd837, 32'sd935,
32'sd915, 32'sd1790, 32'sd501, 32'sd1544, 32'sd226, 32'sd269,
32'sd1799, 32'sd659, 32'sd966, 32'sd1150, 32'sd716, 32'sd1332,
32'sd1547, 32'sd1251, 32'sd1838, 32'sd1644, 32'sd1509, 32'sd1313,
32'sd1997, 32'sd1807, 32'sd1329, 32'sd1957, 32'sd1719, 32'sd620,
32'sd208, 32'sd488, 32'sd642, 32'sd306, 32'sd447, 32'sd693,
32'sd1394, 32'sd552, 32'sd362, 32'sd1617, 32'sd1137, 32'sd820,
32'sd1570, 32'sd537, 32'sd1670, 32'sd1408, 32'sd1724, 32'sd1710,
32'sd1123, 32'sd1351, 32'sd1300, 32'sd141, 32'sd1164, 32'sd1187,
32'sd734, 32'sd743, 32'sd1501, 32'sd1265, 32'sd106, 32'sd1472,
32'sd1064, 32'sd865, 32'sd1403, 32'sd504, 32'sd1518, 32'sd1283,
32'sd352, 32'sd359, 32'sd1833, 32'sd1877, 32'sd465, 32'sd1396,
32'sd170, 32'sd1501, 32'sd602, 32'sd925, 32'sd1373, 32'sd982,
32'sd408, 32'sd747, 32'sd1762, 32'sd406, 32'sd942, 32'sd738,
32'sd323, 32'sd1947, 32'sd1834, 32'sd532, 32'sd380, 32'sd1676,
32'sd1163, 32'sd1631, 32'sd836, 32'sd1434, 32'sd1527, 32'sd1331,
32'sd1639, 32'sd1550, 32'sd1656, 32'sd945, 32'sd1998, 32'sd134,
32'sd372, 32'sd329, 32'sd1697, 32'sd1209, 32'sd802, 32'sd1270,
32'sd1969, 32'sd506, 32'sd423, 32'sd341, 32'sd540, 32'sd255,
32'sd455, 32'sd1232, 32'sd260, 32'sd973, 32'sd1919, 32'sd704,
32'sd1346, 32'sd122, 32'sd453, 32'sd915, 32'sd1865, 32'sd140,
32'sd1422, 32'sd347, 32'sd797, 32'sd231, 32'sd548, 32'sd1687,
32'sd1606, 32'sd1121, 32'sd794, 32'sd1029, 32'sd950, 32'sd170,
32'sd609, 32'sd1694, 32'sd1102, 32'sd1330, 32'sd1071, 32'sd1407,
32'sd1483, 32'sd182, 32'sd228, 32'sd758, 32'sd1733, 32'sd947,
32'sd1067, 32'sd530, 32'sd1198, 32'sd1206, 32'sd767, 32'sd807,
32'sd1451, 32'sd1026, 32'sd1518, 32'sd348, 32'sd1213, 32'sd1470,
32'sd924, 32'sd1336, 32'sd1906, 32'sd783, 32'sd319, 32'sd755,
32'sd1043, 32'sd451, 32'sd974, 32'sd815, 32'sd438, 32'sd1432,
32'sd1464, 32'sd1970, 32'sd1403, 32'sd879, 32'sd339, 32'sd183,
32'sd369, 32'sd765, 32'sd771, 32'sd1958, 32'sd553, 32'sd334,
32'sd825, 32'sd906, 32'sd1323, 32'sd1712, 32'sd979, 32'sd133,
32'sd1951, 32'sd366, 32'sd826, 32'sd798, 32'sd1550, 32'sd513,
32'sd766, 32'sd280, 32'sd299, 32'sd1463, 32'sd1171, 32'sd139,
32'sd191, 32'sd200, 32'sd582, 32'sd1514, 32'sd789, 32'sd1432,
32'sd319, 32'sd1026, 32'sd1911, 32'sd1733, 32'sd329, 32'sd970,
32'sd1043, 32'sd997, 32'sd437, 32'sd1047, 32'sd578, 32'sd1257,
32'sd1188, 32'sd1917, 32'sd1778, 32'sd1508, 32'sd587, 32'sd352,
32'sd534, 32'sd816, 32'sd404, 32'sd625, 32'sd1044, 32'sd1931,
32'sd1654, 32'sd1222, 32'sd1384, 32'sd1905, 32'sd870, 32'sd890,
32'sd1440, 32'sd815, 32'sd552, 32'sd411, 32'sd1319, 32'sd1588,
32'sd278, 32'sd102, 32'sd1413, 32'sd1056, 32'sd1905, 32'sd344,
32'sd1504, 32'sd243, 32'sd196, 32'sd1957, 32'sd461, 32'sd677,
32'sd804, 32'sd1682, 32'sd361, 32'sd127, 32'sd883, 32'sd1579,
32'sd1311, 32'sd929, 32'sd1930, 32'sd1256, 32'sd368, 32'sd458,
32'sd191, 32'sd843, 32'sd1722, 32'sd938, 32'sd107, 32'sd511,
32'sd1472, 32'sd1601, 32'sd1510, 32'sd249, 32'sd1145, 32'sd1309,
32'sd803, 32'sd257, 32'sd1646, 32'sd126, 32'sd1247, 32'sd1072,
32'sd1497, 32'sd463, 32'sd287, 32'sd408, 32'sd399, 32'sd892,
32'sd1272, 32'sd959, 32'sd498, 32'sd293, 32'sd1587, 32'sd582,
32'sd1005, 32'sd1149, 32'sd841, 32'sd1064, 32'sd956, 32'sd1689,
32'sd1212, 32'sd209, 32'sd659, 32'sd1131, 32'sd585, 32'sd1431,
32'sd492, 32'sd341, 32'sd1408, 32'sd1706, 32'sd1933, 32'sd1268,
32'sd293, 32'sd1919, 32'sd1839, 32'sd1326, 32'sd1228, 32'sd920,
32'sd1894, 32'sd1194, 32'sd1039, 32'sd416, 32'sd1953, 32'sd340,
32'sd466, 32'sd1193, 32'sd1484, 32'sd1563, 32'sd473, 32'sd254,
32'sd418, 32'sd201, 32'sd1774, 32'sd788, 32'sd319, 32'sd1191,
32'sd596, 32'sd1189, 32'sd897, 32'sd1489, 32'sd1047, 32'sd594,
32'sd1676, 32'sd530, 32'sd618, 32'sd1071, 32'sd1694, 32'sd1028,
32'sd374, 32'sd217, 32'sd1814, 32'sd1297, 32'sd1845, 32'sd1991,
32'sd1349, 32'sd1947, 32'sd1981, 32'sd1542, 32'sd524, 32'sd1893,
32'sd702, 32'sd933, 32'sd803, 32'sd408, 32'sd1797, 32'sd1195,
32'sd1851, 32'sd1196, 32'sd499, 32'sd445, 32'sd1100, 32'sd948,
32'sd1726, 32'sd1493, 32'sd1230, 32'sd297, 32'sd1987, 32'sd1063,
32'sd311, 32'sd232, 32'sd1500, 32'sd436, 32'sd1067, 32'sd394,
32'sd327, 32'sd184, 32'sd1696, 32'sd767, 32'sd1023, 32'sd1916,
32'sd926, 32'sd1659, 32'sd201, 32'sd802, 32'sd157, 32'sd200,
32'sd194, 32'sd242, 32'sd1770, 32'sd111, 32'sd1598, 32'sd1402,
32'sd564, 32'sd1772, 32'sd1452, 32'sd301, 32'sd1958, 32'sd172,
32'sd590, 32'sd194, 32'sd573, 32'sd1092, 32'sd1025, 32'sd1977,
32'sd441, 32'sd426, 32'sd103, 32'sd653, 32'sd1723, 32'sd1673,
32'sd608, 32'sd1992, 32'sd1893, 32'sd478, 32'sd655, 32'sd1671,
32'sd833, 32'sd1840, 32'sd848, 32'sd1891, 32'sd1085, 32'sd111,
32'sd571, 32'sd441, 32'sd1181, 32'sd724, 32'sd574, 32'sd790,
32'sd413, 32'sd1906, 32'sd1373, 32'sd1645, 32'sd112, 32'sd1872,
32'sd876, 32'sd1548, 32'sd1347, 32'sd844, 32'sd289, 32'sd1336,
32'sd838, 32'sd620, 32'sd747, 32'sd641, 32'sd1001, 32'sd1328,
32'sd201, 32'sd713, 32'sd227, 32'sd857, 32'sd1615, 32'sd1282,
32'sd1245, 32'sd1804, 32'sd442, 32'sd1280, 32'sd1095, 32'sd505,
32'sd944, 32'sd220, 32'sd842, 32'sd1229, 32'sd1112, 32'sd1426,
32'sd397, 32'sd1333, 32'sd338, 32'sd477, 32'sd1504, 32'sd1125,
32'sd833, 32'sd1766, 32'sd1720, 32'sd1485, 32'sd646, 32'sd1550,
32'sd1311, 32'sd1596, 32'sd924, 32'sd1528, 32'sd1842, 32'sd1602,
32'sd345, 32'sd553, 32'sd1260, 32'sd730, 32'sd562, 32'sd1030,
32'sd334, 32'sd1742, 32'sd1079, 32'sd573, 32'sd1332, 32'sd1842,
32'sd181, 32'sd342, 32'sd393, 32'sd724, 32'sd782, 32'sd210,
32'sd237, 32'sd133, 32'sd195, 32'sd405, 32'sd1985, 32'sd1095,
32'sd336, 32'sd1595, 32'sd1005, 32'sd1196, 32'sd1759, 32'sd449,
32'sd1430, 32'sd823, 32'sd427, 32'sd803, 32'sd286, 32'sd159,
32'sd655, 32'sd200, 32'sd609, 32'sd915, 32'sd214, 32'sd201,
32'sd764, 32'sd709, 32'sd1976, 32'sd1115, 32'sd1717, 32'sd1770,
32'sd1587, 32'sd147, 32'sd542, 32'sd1704, 32'sd1859, 32'sd238,
32'sd1397, 32'sd131, 32'sd1135, 32'sd219, 32'sd1743, 32'sd1813,
32'sd670, 32'sd392, 32'sd1137, 32'sd698, 32'sd990, 32'sd303,
32'sd313, 32'sd1979, 32'sd461, 32'sd571, 32'sd1527, 32'sd1958,
32'sd1170, 32'sd209, 32'sd857, 32'sd1308, 32'sd1751, 32'sd1819,
32'sd1098, 32'sd1865, 32'sd1677, 32'sd1060, 32'sd1116, 32'sd623,
32'sd1853, 32'sd451, 32'sd527, 32'sd1174, 32'sd738, 32'sd1839,
32'sd1244, 32'sd1885, 32'sd1134, 32'sd1568, 32'sd1245, 32'sd1714,
32'sd691, 32'sd1709, 32'sd1403, 32'sd270, 32'sd1522, 32'sd1330,
32'sd225, 32'sd597, 32'sd1044, 32'sd1299, 32'sd299, 32'sd1921,
32'sd1508, 32'sd680, 32'sd1818, 32'sd1285, 32'sd1899, 32'sd1182,
32'sd1754, 32'sd698, 32'sd912, 32'sd875, 32'sd1906, 32'sd829,
32'sd932, 32'sd853, 32'sd447, 32'sd1319, 32'sd1363, 32'sd1444,
32'sd888, 32'sd1151, 32'sd791, 32'sd486, 32'sd273, 32'sd396,
32'sd112, 32'sd1588, 32'sd620, 32'sd1932, 32'sd532, 32'sd1300,
32'sd1312, 32'sd788, 32'sd1855, 32'sd524, 32'sd1288, 32'sd1838,
32'sd1933, 32'sd130, 32'sd1263, 32'sd1662, 32'sd838, 32'sd907,
32'sd1404, 32'sd971, 32'sd1234, 32'sd1469, 32'sd1041, 32'sd1509,
32'sd1195, 32'sd1257, 32'sd1648, 32'sd639, 32'sd1487, 32'sd170,
32'sd191, 32'sd1225, 32'sd1446, 32'sd1547, 32'sd193, 32'sd1841,
32'sd714, 32'sd1652, 32'sd1862, 32'sd632, 32'sd1949, 32'sd1584,
32'sd1116, 32'sd1403, 32'sd1866, 32'sd944, 32'sd876, 32'sd1675,
32'sd307, 32'sd1678, 32'sd463, 32'sd1817, 32'sd1577, 32'sd522,
32'sd1953, 32'sd428, 32'sd1404, 32'sd933, 32'sd478, 32'sd1228,
32'sd611, 32'sd426, 32'sd924, 32'sd1027, 32'sd673, 32'sd1593,
32'sd1784, 32'sd201, 32'sd583, 32'sd1470, 32'sd1607, 32'sd1663,
32'sd619, 32'sd1350, 32'sd671, 32'sd1713, 32'sd729, 32'sd1207,
32'sd1994, 32'sd1587, 32'sd1277, 32'sd557, 32'sd250, 32'sd1692,
32'sd1997, 32'sd1889, 32'sd1129, 32'sd152, 32'sd158, 32'sd1668,
32'sd198, 32'sd1047, 32'sd1336, 32'sd1830, 32'sd1246, 32'sd1719,
32'sd1602, 32'sd259, 32'sd1428, 32'sd1865, 32'sd890, 32'sd734,
32'sd812, 32'sd1297, 32'sd1188, 32'sd1412, 32'sd1191, 32'sd1641,
32'sd1061, 32'sd155, 32'sd811, 32'sd1758, 32'sd1669, 32'sd141,
32'sd837, 32'sd207, 32'sd106, 32'sd830, 32'sd529, 32'sd1195,
32'sd679, 32'sd934, 32'sd1021, 32'sd679, 32'sd1877, 32'sd1310,
32'sd1005, 32'sd116, 32'sd155, 32'sd1202, 32'sd1324, 32'sd1518,
32'sd334, 32'sd290, 32'sd1921, 32'sd1976, 32'sd510, 32'sd381,
32'sd1040, 32'sd1339, 32'sd773, 32'sd284, 32'sd1788, 32'sd1320,
32'sd1726, 32'sd762, 32'sd484, 32'sd166, 32'sd802, 32'sd1117,
32'sd369, 32'sd533, 32'sd1411, 32'sd745, 32'sd1376, 32'sd561,
32'sd918, 32'sd1870, 32'sd669, 32'sd1117, 32'sd422, 32'sd1728,
32'sd474, 32'sd1846, 32'sd972, 32'sd684, 32'sd1807, 32'sd1268,
32'sd836, 32'sd1118, 32'sd1623, 32'sd1013, 32'sd415, 32'sd238,
32'sd403, 32'sd1955, 32'sd279, 32'sd271, 32'sd1709, 32'sd436,
32'sd1072, 32'sd1565, 32'sd124, 32'sd1679, 32'sd1426, 32'sd945,
32'sd1976, 32'sd658, 32'sd1588, 32'sd1110, 32'sd1642, 32'sd1655,
32'sd809, 32'sd559, 32'sd1814, 32'sd1775, 32'sd1640, 32'sd1464,
32'sd225, 32'sd1760, 32'sd1712, 32'sd218, 32'sd1710, 32'sd849,
32'sd1172, 32'sd402, 32'sd334, 32'sd395, 32'sd411, 32'sd1904,
32'sd1771, 32'sd128, 32'sd1587, 32'sd449, 32'sd622, 32'sd1868,
32'sd132, 32'sd871, 32'sd543, 32'sd1147, 32'sd908, 32'sd384,
32'sd1762, 32'sd309, 32'sd231, 32'sd1310, 32'sd871, 32'sd1738,
32'sd189, 32'sd1526, 32'sd1853, 32'sd578, 32'sd970, 32'sd1073,
32'sd890, 32'sd568, 32'sd866, 32'sd578, 32'sd1085, 32'sd1384,
32'sd1282, 32'sd1639, 32'sd1427, 32'sd1518, 32'sd1425, 32'sd1470,
32'sd1045, 32'sd887, 32'sd516, 32'sd1461, 32'sd1224, 32'sd239,
32'sd448, 32'sd644, 32'sd1653, 32'sd930, 32'sd460, 32'sd238,
32'sd611, 32'sd1868, 32'sd797, 32'sd823, 32'sd235, 32'sd620,
32'sd1287, 32'sd1306, 32'sd618, 32'sd408, 32'sd465, 32'sd388,
32'sd1336, 32'sd726, 32'sd168, 32'sd1719, 32'sd395, 32'sd379,
32'sd488, 32'sd710, 32'sd1264, 32'sd956, 32'sd1585, 32'sd1318,
32'sd1825, 32'sd1970, 32'sd323, 32'sd174, 32'sd1168, 32'sd1884,
32'sd324, 32'sd1031, 32'sd118, 32'sd1147, 32'sd643, 32'sd1815,
32'sd1077, 32'sd1043, 32'sd1557, 32'sd663, 32'sd933, 32'sd608,
32'sd1325, 32'sd1655, 32'sd915, 32'sd662, 32'sd1890, 32'sd1415,
32'sd329, 32'sd980, 32'sd1690, 32'sd1149, 32'sd150, 32'sd1210,
32'sd316, 32'sd989, 32'sd302, 32'sd1712, 32'sd952, 32'sd1906,
32'sd744, 32'sd1127, 32'sd1334, 32'sd732, 32'sd570, 32'sd1971,
32'sd1692, 32'sd1244, 32'sd1476, 32'sd1892, 32'sd162, 32'sd716,
32'sd1509, 32'sd1286, 32'sd972, 32'sd1493, 32'sd1654, 32'sd1252,
32'sd502, 32'sd292, 32'sd802, 32'sd1069, 32'sd1366, 32'sd1103,
32'sd306, 32'sd1981, 32'sd365, 32'sd490, 32'sd1018, 32'sd1305,
32'sd1259, 32'sd928, 32'sd1023, 32'sd500, 32'sd976, 32'sd551,
32'sd1848, 32'sd352, 32'sd1129, 32'sd1150, 32'sd1461, 32'sd344,
32'sd698, 32'sd458, 32'sd1962, 32'sd636, 32'sd310, 32'sd702,
32'sd1063, 32'sd537, 32'sd503, 32'sd636, 32'sd889, 32'sd1801,
32'sd206, 32'sd691, 32'sd568, 32'sd419, 32'sd551, 32'sd742,
32'sd1675, 32'sd828, 32'sd812, 32'sd1128, 32'sd1333, 32'sd1208,
32'sd881, 32'sd1799, 32'sd1637, 32'sd1726, 32'sd815, 32'sd1182,
32'sd1488, 32'sd1369, 32'sd240, 32'sd919, 32'sd230, 32'sd346,
32'sd1731, 32'sd1528, 32'sd1809, 32'sd643, 32'sd1131, 32'sd1258,
32'sd499, 32'sd1480, 32'sd1353, 32'sd1520, 32'sd1801, 32'sd1743,
32'sd575, 32'sd1688, 32'sd1117, 32'sd704, 32'sd1003, 32'sd334,
32'sd1041, 32'sd1690, 32'sd1698, 32'sd1523, 32'sd378, 32'sd1701,
32'sd1870, 32'sd517, 32'sd1962, 32'sd278, 32'sd169, 32'sd1063,
32'sd709, 32'sd1153, 32'sd1163, 32'sd834, 32'sd809, 32'sd615,
32'sd184, 32'sd1952, 32'sd934, 32'sd1616, 32'sd501, 32'sd1078,
32'sd714, 32'sd194, 32'sd290, 32'sd1146, 32'sd1517, 32'sd1588,
32'sd1138, 32'sd671, 32'sd1802, 32'sd1474, 32'sd224, 32'sd1991,
32'sd1393, 32'sd595, 32'sd1043, 32'sd844, 32'sd1947, 32'sd478,
32'sd886, 32'sd1836, 32'sd1112, 32'sd1737, 32'sd728, 32'sd322,
32'sd442, 32'sd1832, 32'sd437, 32'sd463, 32'sd1352, 32'sd261,
32'sd515, 32'sd1270, 32'sd1610, 32'sd1538, 32'sd265, 32'sd726,
32'sd513, 32'sd1907, 32'sd1521, 32'sd407, 32'sd1736, 32'sd939,
32'sd316, 32'sd240, 32'sd811, 32'sd315, 32'sd771, 32'sd1709,
32'sd1086, 32'sd1639, 32'sd676, 32'sd1278, 32'sd1533, 32'sd1725,
32'sd1596, 32'sd1437, 32'sd211, 32'sd1055, 32'sd1890, 32'sd1070,
32'sd1834, 32'sd1731, 32'sd495, 32'sd569, 32'sd166, 32'sd995,
32'sd674, 32'sd122, 32'sd604, 32'sd134, 32'sd297, 32'sd1855,
32'sd470, 32'sd1402, 32'sd1685, 32'sd621, 32'sd1616, 32'sd493,
32'sd692, 32'sd1139, 32'sd327, 32'sd580, 32'sd1734, 32'sd1418,
32'sd550, 32'sd403, 32'sd783, 32'sd599, 32'sd1392, 32'sd836,
32'sd387, 32'sd1083, 32'sd414, 32'sd1373, 32'sd111, 32'sd1849,
32'sd654, 32'sd1621, 32'sd986, 32'sd889, 32'sd340, 32'sd710,
32'sd1391, 32'sd208, 32'sd419, 32'sd1963, 32'sd1541, 32'sd1793,
32'sd1746, 32'sd329, 32'sd1365, 32'sd760, 32'sd468, 32'sd979,
32'sd262, 32'sd815, 32'sd1636, 32'sd1976, 32'sd1831, 32'sd1435,
32'sd1772, 32'sd924, 32'sd1295, 32'sd1794, 32'sd1711, 32'sd665,
32'sd1966, 32'sd908, 32'sd368, 32'sd1735, 32'sd580, 32'sd1571,
32'sd776, 32'sd805, 32'sd324, 32'sd371, 32'sd1215, 32'sd225,
32'sd1413, 32'sd362, 32'sd691, 32'sd922, 32'sd351, 32'sd245,
32'sd1776, 32'sd1490, 32'sd727, 32'sd782, 32'sd188, 32'sd1994,
32'sd1683, 32'sd1369, 32'sd181, 32'sd1822, 32'sd1620, 32'sd873,
32'sd1337, 32'sd210, 32'sd1727, 32'sd1924, 32'sd954, 32'sd933,
32'sd1373, 32'sd1175, 32'sd974, 32'sd774, 32'sd1230, 32'sd1146,
32'sd559, 32'sd1521, 32'sd452, 32'sd880, 32'sd562, 32'sd161,
32'sd607, 32'sd480, 32'sd1710, 32'sd259, 32'sd1122, 32'sd251,
32'sd1085, 32'sd1624, 32'sd1292, 32'sd225, 32'sd1374, 32'sd1737,
32'sd1858, 32'sd1004, 32'sd1177, 32'sd1786, 32'sd1044, 32'sd1698,
32'sd1716, 32'sd1483, 32'sd1083, 32'sd158, 32'sd1527, 32'sd1961,
32'sd144, 32'sd729, 32'sd1400, 32'sd973, 32'sd1584, 32'sd201,
32'sd1681, 32'sd994, 32'sd1054, 32'sd158, 32'sd1722, 32'sd1887,
32'sd1280, 32'sd771, 32'sd226, 32'sd662, 32'sd1835, 32'sd882,
32'sd470, 32'sd1923, 32'sd503, 32'sd145, 32'sd1080, 32'sd453,
32'sd819, 32'sd226, 32'sd1800, 32'sd441, 32'sd305, 32'sd398,
32'sd1120, 32'sd114, 32'sd1347, 32'sd180, 32'sd1641, 32'sd585,
32'sd548, 32'sd600, 32'sd1001, 32'sd722, 32'sd171, 32'sd239,
32'sd644, 32'sd292, 32'sd1938, 32'sd160, 32'sd1137, 32'sd643,
32'sd481, 32'sd1695, 32'sd1109, 32'sd151, 32'sd1058, 32'sd1893,
32'sd1099, 32'sd1440, 32'sd240, 32'sd916, 32'sd1011, 32'sd822,
32'sd1269, 32'sd721, 32'sd845, 32'sd112, 32'sd855, 32'sd1856,
32'sd892, 32'sd736, 32'sd1967, 32'sd484, 32'sd1968, 32'sd146,
32'sd480, 32'sd869, 32'sd1975, 32'sd141, 32'sd1010, 32'sd619,
32'sd357, 32'sd1711, 32'sd503, 32'sd1990, 32'sd359, 32'sd1749,
32'sd1715, 32'sd329, 32'sd793, 32'sd929, 32'sd1958, 32'sd1478,
32'sd1776, 32'sd1990, 32'sd1791, 32'sd123, 32'sd997, 32'sd216,
32'sd646, 32'sd1968, 32'sd1821, 32'sd812, 32'sd1523, 32'sd539,
32'sd1105, 32'sd1810, 32'sd393, 32'sd1069, 32'sd810, 32'sd1456,
32'sd520, 32'sd542, 32'sd1911, 32'sd688, 32'sd618, 32'sd1708,
32'sd1556, 32'sd313, 32'sd1247, 32'sd1536, 32'sd1782, 32'sd1510,
32'sd1093, 32'sd1121, 32'sd181, 32'sd1182, 32'sd727, 32'sd1272,
32'sd1704, 32'sd1949, 32'sd1016, 32'sd1781, 32'sd1263, 32'sd1294,
32'sd207, 32'sd1814, 32'sd570, 32'sd242, 32'sd1578, 32'sd1907,
32'sd612, 32'sd604, 32'sd766, 32'sd1043, 32'sd1729, 32'sd894,
32'sd151, 32'sd1364, 32'sd993, 32'sd1591, 32'sd1995, 32'sd358,
32'sd187, 32'sd368, 32'sd1192, 32'sd1564, 32'sd738, 32'sd1642,
32'sd456, 32'sd1211, 32'sd1567, 32'sd891, 32'sd974, 32'sd756,
32'sd588, 32'sd1206, 32'sd1807, 32'sd1888, 32'sd1673, 32'sd1258,
32'sd530, 32'sd339, 32'sd1110, 32'sd1948, 32'sd919, 32'sd1272,
32'sd462, 32'sd1001, 32'sd1374, 32'sd1869, 32'sd1222, 32'sd1444,
32'sd821, 32'sd1115, 32'sd214, 32'sd1506, 32'sd1548, 32'sd1479,
32'sd1719, 32'sd880, 32'sd1127, 32'sd189, 32'sd250, 32'sd832,
32'sd401, 32'sd1733, 32'sd1144, 32'sd471, 32'sd1786, 32'sd972,
32'sd1178, 32'sd1047, 32'sd1629, 32'sd190, 32'sd1981, 32'sd549,
32'sd868, 32'sd280, 32'sd1963, 32'sd1874, 32'sd1463, 32'sd713,
32'sd379, 32'sd1713, 32'sd302, 32'sd1320, 32'sd1148, 32'sd1208,
32'sd1201, 32'sd752, 32'sd992, 32'sd707, 32'sd499, 32'sd496,
32'sd1919, 32'sd1927, 32'sd520, 32'sd1652, 32'sd925, 32'sd1573,
32'sd1264, 32'sd1019, 32'sd1988, 32'sd828, 32'sd1771, 32'sd1500,
32'sd513, 32'sd1940, 32'sd324, 32'sd992, 32'sd1817, 32'sd124,
32'sd1153, 32'sd1546, 32'sd1411, 32'sd930, 32'sd1006, 32'sd1227,
32'sd1641, 32'sd491, 32'sd578, 32'sd1471, 32'sd1832, 32'sd1987,
32'sd329, 32'sd537, 32'sd1265, 32'sd201, 32'sd1363, 32'sd862,
32'sd462, 32'sd1950, 32'sd1016, 32'sd805, 32'sd1884, 32'sd309,
32'sd1492, 32'sd350, 32'sd990, 32'sd1645, 32'sd580, 32'sd235,
32'sd1183, 32'sd1460, 32'sd592, 32'sd1243, 32'sd1288, 32'sd1783,
32'sd597, 32'sd294, 32'sd1532, 32'sd1172, 32'sd1637, 32'sd415,
32'sd206, 32'sd1536, 32'sd1530, 32'sd134, 32'sd1222, 32'sd724,
32'sd1065, 32'sd1292, 32'sd1855, 32'sd586, 32'sd228, 32'sd157,
32'sd1366, 32'sd632, 32'sd1689, 32'sd1348, 32'sd1097, 32'sd490,
32'sd1795, 32'sd1366, 32'sd1176, 32'sd268, 32'sd333, 32'sd1722,
32'sd336, 32'sd382, 32'sd741, 32'sd1116, 32'sd531, 32'sd990,
32'sd215, 32'sd876, 32'sd1465, 32'sd1769, 32'sd1812, 32'sd1484,
32'sd1963, 32'sd1220, 32'sd552, 32'sd1564, 32'sd1073, 32'sd1280,
32'sd1957, 32'sd682, 32'sd840, 32'sd888, 32'sd1160, 32'sd1099,
32'sd1099, 32'sd974, 32'sd620, 32'sd1971, 32'sd1807, 32'sd511,
32'sd254, 32'sd321, 32'sd1706, 32'sd1028, 32'sd1856, 32'sd200,
32'sd1724, 32'sd1054, 32'sd706, 32'sd720, 32'sd1730, 32'sd789,
32'sd567, 32'sd661, 32'sd880, 32'sd934, 32'sd756, 32'sd1253,
32'sd1487, 32'sd1543, 32'sd544, 32'sd846, 32'sd1976, 32'sd1514,
32'sd1502, 32'sd886, 32'sd362, 32'sd910, 32'sd1804, 32'sd1228,
32'sd1879, 32'sd1232, 32'sd1088, 32'sd1581, 32'sd166, 32'sd937,
32'sd525, 32'sd1673, 32'sd1797, 32'sd1572, 32'sd1156, 32'sd1017,
32'sd1213, 32'sd730, 32'sd1425, 32'sd160, 32'sd1932, 32'sd1010,
32'sd1808, 32'sd1378, 32'sd282, 32'sd1859, 32'sd1275, 32'sd1456,
32'sd194, 32'sd583, 32'sd694, 32'sd358, 32'sd905, 32'sd1671,
32'sd1742, 32'sd1913, 32'sd531, 32'sd458, 32'sd1574, 32'sd1246,
32'sd739, 32'sd1700, 32'sd866, 32'sd941, 32'sd1864, 32'sd1205,
32'sd791, 32'sd1178, 32'sd133, 32'sd1298, 32'sd203, 32'sd441,
32'sd1702, 32'sd298, 32'sd1042, 32'sd438, 32'sd1189, 32'sd879,
32'sd713, 32'sd692, 32'sd866, 32'sd419, 32'sd1425, 32'sd729,
32'sd258, 32'sd338, 32'sd519, 32'sd533, 32'sd1676, 32'sd432,
32'sd899, 32'sd587, 32'sd1546, 32'sd1479, 32'sd670, 32'sd628,
32'sd1682, 32'sd1326, 32'sd170, 32'sd780, 32'sd748, 32'sd357,
32'sd267, 32'sd881, 32'sd1636, 32'sd1048, 32'sd700, 32'sd725,
32'sd1403, 32'sd288, 32'sd1623, 32'sd906, 32'sd584, 32'sd353,
32'sd364, 32'sd993, 32'sd471, 32'sd1178, 32'sd127, 32'sd1776,
32'sd1684, 32'sd700, 32'sd819, 32'sd1725, 32'sd440, 32'sd362,
32'sd1134, 32'sd218, 32'sd1774, 32'sd1906, 32'sd1110, 32'sd1775,
32'sd788, 32'sd264, 32'sd1587, 32'sd1800, 32'sd960, 32'sd581,
32'sd1961, 32'sd370, 32'sd750, 32'sd1829, 32'sd958, 32'sd384,
32'sd1008, 32'sd547, 32'sd1882, 32'sd557, 32'sd890, 32'sd348,
32'sd997, 32'sd1007, 32'sd789, 32'sd1070, 32'sd113, 32'sd1145,
32'sd1545, 32'sd1643, 32'sd376, 32'sd774, 32'sd806, 32'sd1216,
32'sd332, 32'sd1124, 32'sd1687, 32'sd121, 32'sd779, 32'sd1061,
32'sd165, 32'sd1666, 32'sd744, 32'sd1823, 32'sd1722, 32'sd101,
32'sd464, 32'sd346, 32'sd552, 32'sd256, 32'sd1249, 32'sd1196,
32'sd611, 32'sd1294, 32'sd966, 32'sd846, 32'sd116, 32'sd216,
32'sd852, 32'sd1452, 32'sd955, 32'sd1033, 32'sd270, 32'sd1553,
32'sd1307, 32'sd1278, 32'sd1593, 32'sd1309, 32'sd1028, 32'sd1431,
32'sd955, 32'sd981, 32'sd1803, 32'sd504, 32'sd263, 32'sd1297,
32'sd804, 32'sd895, 32'sd1884, 32'sd403, 32'sd1432, 32'sd1136,
32'sd427, 32'sd1455, 32'sd1725, 32'sd377, 32'sd1913, 32'sd1041,
32'sd1564, 32'sd136, 32'sd172, 32'sd731, 32'sd1178, 32'sd585,
32'sd926, 32'sd1679, 32'sd528, 32'sd758, 32'sd943, 32'sd685,
32'sd382, 32'sd1171, 32'sd1967, 32'sd1342, 32'sd1342, 32'sd1199,
32'sd1164, 32'sd1493, 32'sd1001, 32'sd1170, 32'sd159, 32'sd1262,
32'sd1476, 32'sd328, 32'sd226, 32'sd246, 32'sd703, 32'sd547,
32'sd787, 32'sd704, 32'sd262, 32'sd1357, 32'sd1638, 32'sd333,
32'sd1419, 32'sd122, 32'sd1175, 32'sd1402, 32'sd1497, 32'sd1613,
32'sd1002, 32'sd1440, 32'sd907, 32'sd1760, 32'sd1846, 32'sd919,
32'sd1508, 32'sd429, 32'sd985, 32'sd836, 32'sd1352, 32'sd736,
32'sd1167, 32'sd678, 32'sd1111, 32'sd1112, 32'sd1925, 32'sd1632,
32'sd1317, 32'sd1542, 32'sd330, 32'sd413, 32'sd1414, 32'sd823,
32'sd1602, 32'sd1309, 32'sd1380, 32'sd1008, 32'sd991, 32'sd1230,
32'sd294, 32'sd1387, 32'sd1894, 32'sd1931, 32'sd1286, 32'sd1082,
32'sd1799, 32'sd546, 32'sd976, 32'sd1274, 32'sd613, 32'sd1175,
32'sd1645, 32'sd102, 32'sd909, 32'sd135, 32'sd503, 32'sd178,
32'sd377, 32'sd527, 32'sd1945, 32'sd1770, 32'sd519, 32'sd1733,
32'sd1540, 32'sd438, 32'sd660, 32'sd1864, 32'sd1843, 32'sd1861,
32'sd951, 32'sd1964, 32'sd880, 32'sd1454, 32'sd356, 32'sd715,
32'sd1821, 32'sd1572, 32'sd199, 32'sd1942, 32'sd706, 32'sd578,
32'sd406, 32'sd507, 32'sd1817, 32'sd1221, 32'sd1383, 32'sd271,
32'sd374, 32'sd538, 32'sd1677, 32'sd520, 32'sd1161, 32'sd994,
32'sd775, 32'sd869, 32'sd1012, 32'sd1536, 32'sd503, 32'sd563,
32'sd496, 32'sd1853, 32'sd110, 32'sd1122, 32'sd1823, 32'sd1594,
32'sd1047, 32'sd1924, 32'sd118, 32'sd1465, 32'sd1873, 32'sd1169,
32'sd583, 32'sd1077, 32'sd1142, 32'sd1962, 32'sd662, 32'sd931,
32'sd1631, 32'sd681, 32'sd1472, 32'sd813, 32'sd660, 32'sd1777,
32'sd150, 32'sd880, 32'sd826, 32'sd144, 32'sd1189, 32'sd1278,
32'sd1852, 32'sd800, 32'sd1176, 32'sd1951, 32'sd1832, 32'sd871,
32'sd976, 32'sd1055, 32'sd353, 32'sd290, 32'sd1294, 32'sd1270,
32'sd645, 32'sd1785, 32'sd426, 32'sd1801, 32'sd215, 32'sd341,
32'sd791, 32'sd261, 32'sd603, 32'sd1719, 32'sd1654, 32'sd390,
32'sd267, 32'sd1522, 32'sd553, 32'sd662, 32'sd1940, 32'sd1156,
32'sd1154, 32'sd1897, 32'sd807, 32'sd803, 32'sd401, 32'sd538,
32'sd206, 32'sd1779, 32'sd1788, 32'sd149, 32'sd1733, 32'sd1204,
32'sd1492, 32'sd1069, 32'sd654, 32'sd749, 32'sd551, 32'sd396,
32'sd737, 32'sd1350, 32'sd1603, 32'sd1646, 32'sd939, 32'sd1385,
32'sd1392, 32'sd1701, 32'sd696, 32'sd1988, 32'sd1183, 32'sd846,
32'sd1249, 32'sd387, 32'sd1517, 32'sd1643, 32'sd967, 32'sd1648,
32'sd1166, 32'sd1344, 32'sd1921, 32'sd550, 32'sd330, 32'sd599,
32'sd934, 32'sd1139, 32'sd1313, 32'sd1792, 32'sd300, 32'sd480,
32'sd1370, 32'sd347, 32'sd1501, 32'sd543, 32'sd1886, 32'sd678,
32'sd1958, 32'sd283, 32'sd777, 32'sd859, 32'sd857, 32'sd162,
32'sd899, 32'sd395, 32'sd1116, 32'sd597, 32'sd118, 32'sd1841,
32'sd1499, 32'sd1721, 32'sd773, 32'sd1447, 32'sd987, 32'sd375,
32'sd960, 32'sd1970, 32'sd741, 32'sd381, 32'sd825, 32'sd1484,
32'sd1866, 32'sd1832, 32'sd114, 32'sd784, 32'sd1993, 32'sd1852,
32'sd1134, 32'sd588, 32'sd584, 32'sd111, 32'sd1041, 32'sd1138,
32'sd1849, 32'sd131, 32'sd680, 32'sd1890, 32'sd1549, 32'sd1947,
32'sd109, 32'sd344, 32'sd985, 32'sd312, 32'sd649, 32'sd1679,
32'sd1593, 32'sd445, 32'sd181, 32'sd788, 32'sd1690, 32'sd1317,
32'sd1131, 32'sd255, 32'sd717, 32'sd1341, 32'sd276, 32'sd290,
32'sd1900, 32'sd995, 32'sd142, 32'sd233, 32'sd1358, 32'sd1790,
32'sd1961, 32'sd1651, 32'sd794, 32'sd266, 32'sd1491, 32'sd173,
32'sd1848, 32'sd784, 32'sd1693, 32'sd1366, 32'sd1968, 32'sd421,
32'sd1655, 32'sd1896, 32'sd1251, 32'sd1253, 32'sd450, 32'sd489,
32'sd890, 32'sd511, 32'sd677, 32'sd1377, 32'sd874, 32'sd217,
32'sd908, 32'sd1188, 32'sd105, 32'sd1800, 32'sd379, 32'sd1028,
32'sd1364, 32'sd1410, 32'sd1124, 32'sd1750, 32'sd992, 32'sd1327,
32'sd1617, 32'sd1833, 32'sd1268, 32'sd1628, 32'sd120, 32'sd1085,
32'sd1832, 32'sd663, 32'sd170, 32'sd188, 32'sd1677, 32'sd834,
32'sd1527, 32'sd1699, 32'sd591, 32'sd1407, 32'sd1560, 32'sd1599,
32'sd590, 32'sd1061, 32'sd1333, 32'sd184, 32'sd352, 32'sd237,
32'sd1140, 32'sd834, 32'sd1466, 32'sd1794, 32'sd1094, 32'sd1874,
32'sd198, 32'sd726, 32'sd1522, 32'sd1849, 32'sd1681, 32'sd383,
32'sd1448, 32'sd1189, 32'sd1797, 32'sd310, 32'sd1599, 32'sd849,
32'sd690, 32'sd1117, 32'sd1677, 32'sd194, 32'sd1571, 32'sd953,
32'sd1290, 32'sd1327, 32'sd1450, 32'sd1164, 32'sd1814, 32'sd1422,
32'sd1392, 32'sd1427, 32'sd843, 32'sd1438, 32'sd1396, 32'sd1905,
32'sd139, 32'sd1445, 32'sd358, 32'sd978, 32'sd1190, 32'sd1917,
32'sd858, 32'sd1536, 32'sd1363, 32'sd273, 32'sd1885, 32'sd407,
32'sd689, 32'sd1411, 32'sd1926, 32'sd1676, 32'sd1117, 32'sd1217,
32'sd943, 32'sd1733, 32'sd1517, 32'sd836, 32'sd1332, 32'sd1511,
32'sd1803, 32'sd492, 32'sd1675, 32'sd602, 32'sd393, 32'sd1645,
32'sd1180, 32'sd420, 32'sd555, 32'sd156, 32'sd1330, 32'sd973,
32'sd1604, 32'sd810, 32'sd1726, 32'sd330, 32'sd232, 32'sd738,
32'sd1807, 32'sd429, 32'sd1007, 32'sd1281, 32'sd875, 32'sd514,
32'sd879, 32'sd318, 32'sd1842, 32'sd1979, 32'sd1876, 32'sd683,
32'sd1895, 32'sd1302, 32'sd1735, 32'sd1914, 32'sd428, 32'sd754,
32'sd905, 32'sd541, 32'sd1906, 32'sd706, 32'sd1833, 32'sd1514,
32'sd1471, 32'sd718, 32'sd1166, 32'sd1880, 32'sd1822, 32'sd1742,
32'sd851, 32'sd1897, 32'sd1036, 32'sd225, 32'sd1859, 32'sd1230,
32'sd1923, 32'sd1391, 32'sd1720, 32'sd360, 32'sd1111, 32'sd599,
32'sd1664, 32'sd739, 32'sd1970, 32'sd1383, 32'sd1670, 32'sd1631,
32'sd1537, 32'sd1456, 32'sd364, 32'sd568, 32'sd316, 32'sd1470,
32'sd968, 32'sd719, 32'sd1768, 32'sd588, 32'sd1760, 32'sd1094,
32'sd150, 32'sd1114, 32'sd343, 32'sd480, 32'sd1809, 32'sd173,
32'sd200, 32'sd1009, 32'sd937, 32'sd112, 32'sd467, 32'sd1091,
32'sd1619, 32'sd1192, 32'sd353, 32'sd196, 32'sd1440, 32'sd1501,
32'sd1091, 32'sd142, 32'sd537, 32'sd1719, 32'sd1352, 32'sd1653,
32'sd183, 32'sd1360, 32'sd1552, 32'sd876, 32'sd476, 32'sd1938,
32'sd645, 32'sd1837, 32'sd169, 32'sd752, 32'sd942, 32'sd760,
32'sd1532, 32'sd877, 32'sd397, 32'sd879, 32'sd1446, 32'sd323,
32'sd1318, 32'sd559, 32'sd1526, 32'sd558, 32'sd1036, 32'sd1582,
32'sd1951, 32'sd1281, 32'sd1697, 32'sd958, 32'sd868, 32'sd648,
32'sd860, 32'sd1908, 32'sd607, 32'sd341, 32'sd594, 32'sd939,
32'sd1628, 32'sd1561, 32'sd887, 32'sd736, 32'sd1802, 32'sd815,
32'sd426, 32'sd1408, 32'sd1043, 32'sd396, 32'sd1917, 32'sd868,
32'sd330, 32'sd1889, 32'sd559, 32'sd500, 32'sd629, 32'sd120,
32'sd757, 32'sd746, 32'sd1110, 32'sd1135, 32'sd223, 32'sd1360,
32'sd1109, 32'sd1748, 32'sd896, 32'sd867, 32'sd1704, 32'sd710,
32'sd665, 32'sd755, 32'sd561, 32'sd678, 32'sd287, 32'sd764,
32'sd538, 32'sd1953, 32'sd1000, 32'sd1664, 32'sd558, 32'sd1182,
32'sd800, 32'sd374, 32'sd1206, 32'sd693, 32'sd605, 32'sd184,
32'sd953, 32'sd638, 32'sd841, 32'sd430, 32'sd141, 32'sd645,
32'sd797, 32'sd853, 32'sd1808, 32'sd133, 32'sd1095, 32'sd1662,
32'sd1820, 32'sd1664, 32'sd829, 32'sd255, 32'sd1624, 32'sd889,
32'sd1425, 32'sd1194, 32'sd1495, 32'sd868, 32'sd1005, 32'sd630,
32'sd1523, 32'sd1287, 32'sd1964, 32'sd807, 32'sd812, 32'sd555,
32'sd109, 32'sd945, 32'sd837, 32'sd630, 32'sd981, 32'sd514,
32'sd993, 32'sd1509, 32'sd709, 32'sd1172, 32'sd1278, 32'sd709,
32'sd1481, 32'sd1896, 32'sd819, 32'sd1173, 32'sd1570, 32'sd185,
32'sd1870, 32'sd1773, 32'sd186, 32'sd1714, 32'sd809, 32'sd1868,
32'sd1565, 32'sd168, 32'sd1566, 32'sd1981, 32'sd1152, 32'sd1471,
32'sd1774, 32'sd1111, 32'sd1077, 32'sd329, 32'sd158, 32'sd1029,
32'sd1809, 32'sd1665, 32'sd560, 32'sd782, 32'sd282, 32'sd238,
32'sd1505, 32'sd1116, 32'sd1174, 32'sd1760, 32'sd563, 32'sd1365,
32'sd103, 32'sd1851, 32'sd1306, 32'sd1275, 32'sd1006, 32'sd328,
32'sd442, 32'sd1503, 32'sd969, 32'sd420, 32'sd1562, 32'sd941,
32'sd1272, 32'sd678, 32'sd959, 32'sd1256, 32'sd1488, 32'sd407,
32'sd1295, 32'sd1978, 32'sd1854, 32'sd506, 32'sd659, 32'sd781,
32'sd1693, 32'sd1561, 32'sd1956, 32'sd1481, 32'sd454, 32'sd488,
32'sd1167, 32'sd1833, 32'sd334, 32'sd348, 32'sd1509, 32'sd1784,
32'sd128, 32'sd105, 32'sd1592, 32'sd531, 32'sd1771, 32'sd668,
32'sd1690, 32'sd736, 32'sd609, 32'sd538, 32'sd241, 32'sd1237,
32'sd1795, 32'sd689, 32'sd475, 32'sd1152, 32'sd1281, 32'sd321,
32'sd1774, 32'sd540, 32'sd1028, 32'sd1034, 32'sd1607, 32'sd1343,
32'sd1497, 32'sd1945, 32'sd1713, 32'sd978, 32'sd1316, 32'sd422,
32'sd1664, 32'sd931, 32'sd1907, 32'sd1241, 32'sd250, 32'sd984,
32'sd1882, 32'sd1251, 32'sd359, 32'sd460, 32'sd1285, 32'sd419,
32'sd718, 32'sd1190, 32'sd181, 32'sd576, 32'sd1880, 32'sd1045,
32'sd1295, 32'sd941, 32'sd1939, 32'sd364, 32'sd291, 32'sd681,
32'sd1591, 32'sd462, 32'sd752, 32'sd1258, 32'sd1184, 32'sd717,
32'sd1627, 32'sd820, 32'sd617, 32'sd1422, 32'sd865, 32'sd657,
32'sd379, 32'sd662, 32'sd1489, 32'sd312, 32'sd1356, 32'sd357,
32'sd1093, 32'sd1373, 32'sd833, 32'sd662, 32'sd186, 32'sd604,
32'sd550, 32'sd602, 32'sd1624, 32'sd345, 32'sd398, 32'sd1742,
32'sd1789, 32'sd618, 32'sd657, 32'sd1977, 32'sd1222, 32'sd1848,
32'sd990, 32'sd861, 32'sd517, 32'sd1514, 32'sd382, 32'sd1075,
32'sd185, 32'sd434, 32'sd1947, 32'sd604, 32'sd1506, 32'sd281,
32'sd954, 32'sd1173, 32'sd1173, 32'sd876, 32'sd686, 32'sd1782,
32'sd327, 32'sd1004, 32'sd1948, 32'sd1862, 32'sd1571, 32'sd927,
32'sd1153, 32'sd951, 32'sd982, 32'sd1614, 32'sd565, 32'sd912,
32'sd465, 32'sd907, 32'sd1961, 32'sd393, 32'sd1597, 32'sd822,
32'sd1349, 32'sd1666, 32'sd1947, 32'sd571, 32'sd868, 32'sd209,
32'sd605, 32'sd730, 32'sd1898, 32'sd238, 32'sd819, 32'sd1206,
32'sd1760, 32'sd1541, 32'sd701, 32'sd1950, 32'sd1786, 32'sd1264,
32'sd682, 32'sd816, 32'sd983, 32'sd1048, 32'sd420, 32'sd1763,
32'sd1009, 32'sd637, 32'sd1482, 32'sd1412, 32'sd1190, 32'sd1864,
32'sd405, 32'sd1228, 32'sd382, 32'sd1669, 32'sd128, 32'sd647,
32'sd568, 32'sd652, 32'sd256, 32'sd1119, 32'sd1363, 32'sd382,
32'sd1946, 32'sd1341, 32'sd1041, 32'sd1476, 32'sd566, 32'sd707,
32'sd595, 32'sd1509, 32'sd951, 32'sd1296, 32'sd488, 32'sd281,
32'sd756, 32'sd945, 32'sd1363, 32'sd1699, 32'sd301, 32'sd1779,
32'sd166, 32'sd1902, 32'sd300, 32'sd212, 32'sd1954, 32'sd449,
32'sd1039, 32'sd1311, 32'sd964, 32'sd1145, 32'sd1674, 32'sd200,
32'sd657, 32'sd1853, 32'sd842, 32'sd1013, 32'sd1353, 32'sd1642,
32'sd1781, 32'sd1991, 32'sd850, 32'sd384, 32'sd623, 32'sd1987,
32'sd563, 32'sd157, 32'sd784, 32'sd843, 32'sd1812, 32'sd1192,
32'sd1847, 32'sd480, 32'sd1426, 32'sd1764, 32'sd420, 32'sd1276,
32'sd374, 32'sd335, 32'sd1114, 32'sd1953, 32'sd1022, 32'sd1020,
32'sd742, 32'sd472, 32'sd1209, 32'sd1173, 32'sd799, 32'sd966,
32'sd1424, 32'sd1016, 32'sd1076, 32'sd1510, 32'sd569, 32'sd1168,
32'sd1313, 32'sd824, 32'sd1776, 32'sd647, 32'sd458, 32'sd1702,
32'sd330, 32'sd174, 32'sd1296, 32'sd1340, 32'sd418, 32'sd593,
32'sd551, 32'sd1854, 32'sd1825, 32'sd255, 32'sd421, 32'sd398,
32'sd1070, 32'sd1786, 32'sd1979, 32'sd388, 32'sd928, 32'sd1235,
32'sd1313, 32'sd901, 32'sd972, 32'sd233, 32'sd1777, 32'sd1898,
32'sd1557, 32'sd1385, 32'sd908, 32'sd117, 32'sd1661, 32'sd444,
32'sd1201, 32'sd1683, 32'sd455, 32'sd1522, 32'sd219, 32'sd1933,
32'sd1436, 32'sd1727, 32'sd1370, 32'sd1667, 32'sd1891, 32'sd1162,
32'sd1667, 32'sd1913, 32'sd489, 32'sd1527, 32'sd236, 32'sd1779,
32'sd1013, 32'sd1675, 32'sd444, 32'sd1405, 32'sd600, 32'sd1145,
32'sd240, 32'sd1697, 32'sd1660, 32'sd1723, 32'sd319, 32'sd1257,
32'sd391, 32'sd1996, 32'sd765, 32'sd1811, 32'sd919, 32'sd733,
32'sd1730, 32'sd902, 32'sd1056, 32'sd348, 32'sd153, 32'sd353,
32'sd1974, 32'sd1056, 32'sd326, 32'sd207, 32'sd162, 32'sd1109,
32'sd1252, 32'sd656, 32'sd1724, 32'sd1291, 32'sd1459, 32'sd1610,
32'sd457, 32'sd148, 32'sd1021, 32'sd394, 32'sd1124, 32'sd193,
32'sd1000, 32'sd1471, 32'sd1253, 32'sd655, 32'sd365, 32'sd933,
32'sd938, 32'sd400, 32'sd570, 32'sd1678, 32'sd983, 32'sd1119,
32'sd1469, 32'sd1646, 32'sd1203, 32'sd1913, 32'sd792, 32'sd130,
32'sd1443, 32'sd398, 32'sd1625, 32'sd103, 32'sd1306, 32'sd1279,
32'sd530, 32'sd1834, 32'sd1667, 32'sd334, 32'sd1793, 32'sd427,
32'sd1833, 32'sd1179, 32'sd930, 32'sd888, 32'sd255, 32'sd1633,
32'sd1520, 32'sd1103, 32'sd605, 32'sd119, 32'sd1042, 32'sd724,
32'sd1563, 32'sd1655, 32'sd1522, 32'sd1475, 32'sd763, 32'sd150,
32'sd527, 32'sd174, 32'sd1630, 32'sd1149, 32'sd1198, 32'sd1786,
32'sd628, 32'sd824, 32'sd467, 32'sd1472, 32'sd1547, 32'sd1341,
32'sd1128, 32'sd1033, 32'sd1334, 32'sd227, 32'sd1463, 32'sd754,
32'sd1830, 32'sd1411, 32'sd665, 32'sd373, 32'sd265, 32'sd1110,
32'sd531, 32'sd1629, 32'sd1010, 32'sd138, 32'sd1607, 32'sd1253,
32'sd952, 32'sd1451, 32'sd346, 32'sd1038, 32'sd1469, 32'sd386,
32'sd524, 32'sd1890, 32'sd1804, 32'sd1289, 32'sd864, 32'sd395,
32'sd1108, 32'sd1411, 32'sd279, 32'sd368, 32'sd1060, 32'sd613,
32'sd1847, 32'sd594, 32'sd1117, 32'sd1636, 32'sd613, 32'sd1833,
32'sd1624, 32'sd235, 32'sd1897, 32'sd1268, 32'sd757, 32'sd1911,
32'sd670, 32'sd833, 32'sd1858, 32'sd1449, 32'sd1808, 32'sd619,
32'sd1284, 32'sd389, 32'sd1012, 32'sd1303, 32'sd1179, 32'sd736,
32'sd479, 32'sd1641, 32'sd251, 32'sd1779, 32'sd1158, 32'sd497,
32'sd1401, 32'sd589, 32'sd568, 32'sd1411, 32'sd1863, 32'sd1100,
32'sd1840, 32'sd1174, 32'sd1325, 32'sd532, 32'sd1698, 32'sd711,
32'sd149, 32'sd1737, 32'sd1609, 32'sd892, 32'sd1783, 32'sd466,
32'sd1979, 32'sd1634, 32'sd1614, 32'sd1286, 32'sd1553, 32'sd1366,
32'sd295, 32'sd891, 32'sd1490, 32'sd1017, 32'sd1547, 32'sd713,
32'sd1299, 32'sd950, 32'sd1331, 32'sd939, 32'sd891, 32'sd1458,
32'sd1068, 32'sd916, 32'sd950, 32'sd310, 32'sd1637, 32'sd385,
32'sd1866, 32'sd496, 32'sd1551, 32'sd1345, 32'sd1859, 32'sd1005,
32'sd274, 32'sd224, 32'sd224, 32'sd1426, 32'sd1446, 32'sd930,
32'sd680, 32'sd572, 32'sd1069, 32'sd1161, 32'sd410, 32'sd927,
32'sd499, 32'sd327, 32'sd1584, 32'sd1687, 32'sd1090, 32'sd1781,
32'sd1996, 32'sd129, 32'sd1474, 32'sd1439, 32'sd497, 32'sd1405,
32'sd639, 32'sd660, 32'sd1494, 32'sd893, 32'sd710, 32'sd412,
32'sd955, 32'sd1696, 32'sd1245, 32'sd257, 32'sd1147, 32'sd1863,
32'sd711, 32'sd1980, 32'sd1701, 32'sd818, 32'sd1630, 32'sd1472,
32'sd1441, 32'sd399, 32'sd572, 32'sd583, 32'sd547, 32'sd648,
32'sd1781, 32'sd584, 32'sd1704, 32'sd1452, 32'sd1936, 32'sd708,
32'sd293, 32'sd702, 32'sd1445, 32'sd470, 32'sd1493, 32'sd564,
32'sd872, 32'sd1923, 32'sd1811, 32'sd771, 32'sd745, 32'sd361,
32'sd1576, 32'sd1370, 32'sd1751, 32'sd1706, 32'sd340, 32'sd737,
32'sd856, 32'sd1778, 32'sd648, 32'sd375, 32'sd538, 32'sd265,
32'sd1326, 32'sd1531, 32'sd455, 32'sd720, 32'sd193, 32'sd1486,
32'sd122, 32'sd1303, 32'sd111, 32'sd1008, 32'sd673, 32'sd1534,
32'sd462, 32'sd1015, 32'sd1648, 32'sd265, 32'sd1361, 32'sd934,
32'sd1623, 32'sd152, 32'sd740, 32'sd141, 32'sd806, 32'sd294,
32'sd1965, 32'sd1906, 32'sd437, 32'sd724, 32'sd1728, 32'sd134,
32'sd1923, 32'sd401, 32'sd947, 32'sd1797, 32'sd1385, 32'sd1386,
32'sd1409, 32'sd1817, 32'sd584, 32'sd1522, 32'sd288, 32'sd1156,
32'sd699, 32'sd1312, 32'sd1979, 32'sd818, 32'sd1736, 32'sd1374,
32'sd1154, 32'sd338, 32'sd1697, 32'sd434, 32'sd496, 32'sd1339,
32'sd1443, 32'sd537, 32'sd709, 32'sd1680, 32'sd1433, 32'sd1339,
32'sd918, 32'sd1209, 32'sd1521, 32'sd494, 32'sd539, 32'sd956,
32'sd926, 32'sd1534, 32'sd725, 32'sd1996, 32'sd1830, 32'sd1854,
32'sd1779, 32'sd808, 32'sd1754, 32'sd128, 32'sd291, 32'sd949,
32'sd1661, 32'sd898, 32'sd1938, 32'sd248, 32'sd1019, 32'sd269,
32'sd436, 32'sd645, 32'sd1409, 32'sd1432, 32'sd874, 32'sd1952,
32'sd1100, 32'sd1142, 32'sd1631, 32'sd684, 32'sd1699, 32'sd1883,
32'sd1838, 32'sd789, 32'sd977, 32'sd655, 32'sd1444, 32'sd743,
32'sd378, 32'sd1914, 32'sd1887, 32'sd244, 32'sd1780, 32'sd1791,
32'sd1818, 32'sd731, 32'sd750, 32'sd152, 32'sd1919, 32'sd1153,
32'sd603, 32'sd576, 32'sd1875, 32'sd607, 32'sd1406, 32'sd1133,
32'sd602, 32'sd1834, 32'sd226, 32'sd1767, 32'sd1073, 32'sd1079,
32'sd219, 32'sd562, 32'sd781, 32'sd294, 32'sd1936, 32'sd1067,
32'sd1155, 32'sd177, 32'sd289, 32'sd500, 32'sd709, 32'sd1825,
32'sd1502, 32'sd419, 32'sd1894, 32'sd283, 32'sd431, 32'sd1147,
32'sd1856, 32'sd1577, 32'sd230, 32'sd1936, 32'sd992, 32'sd1339,
32'sd1744, 32'sd780, 32'sd1631, 32'sd1681, 32'sd1572, 32'sd325,
32'sd1289, 32'sd573, 32'sd1612, 32'sd1946, 32'sd468, 32'sd1632,
32'sd1795, 32'sd1496, 32'sd490, 32'sd291, 32'sd436, 32'sd754,
32'sd168, 32'sd767, 32'sd1877, 32'sd380, 32'sd399, 32'sd1448,
32'sd1118, 32'sd139, 32'sd977, 32'sd600, 32'sd1826, 32'sd309,
32'sd284, 32'sd666, 32'sd1849, 32'sd197, 32'sd1905, 32'sd1507,
32'sd365, 32'sd454, 32'sd172, 32'sd1982, 32'sd1826, 32'sd1040,
32'sd1857, 32'sd1136, 32'sd645, 32'sd1391, 32'sd1349, 32'sd1759,
32'sd1401, 32'sd1894, 32'sd287, 32'sd211, 32'sd684, 32'sd986,
32'sd1120, 32'sd278, 32'sd1911, 32'sd1924, 32'sd735, 32'sd1468,
32'sd105, 32'sd366, 32'sd1636, 32'sd1492, 32'sd1304, 32'sd381,
32'sd827, 32'sd1537, 32'sd1983, 32'sd1616, 32'sd513, 32'sd262,
32'sd779, 32'sd1950, 32'sd466, 32'sd150, 32'sd732, 32'sd831,
32'sd579, 32'sd1963, 32'sd1463, 32'sd1733, 32'sd1750, 32'sd506,
32'sd1704, 32'sd919, 32'sd1134, 32'sd611, 32'sd222, 32'sd380,
32'sd1102, 32'sd1520, 32'sd1487, 32'sd1754, 32'sd688, 32'sd665,
32'sd315, 32'sd1979, 32'sd1330, 32'sd1123, 32'sd823, 32'sd1837,
32'sd1766, 32'sd163, 32'sd282, 32'sd1746, 32'sd1192, 32'sd157,
32'sd1298, 32'sd1275, 32'sd395, 32'sd1697, 32'sd1920, 32'sd168,
32'sd1975, 32'sd1537, 32'sd901, 32'sd510, 32'sd806, 32'sd781,
32'sd1050, 32'sd1519, 32'sd622, 32'sd951, 32'sd1191, 32'sd1096,
32'sd630, 32'sd325, 32'sd1851, 32'sd610, 32'sd991, 32'sd1531,
32'sd1347, 32'sd1369, 32'sd1001, 32'sd1505, 32'sd1220, 32'sd1350,
32'sd727, 32'sd891, 32'sd657, 32'sd1345, 32'sd1097, 32'sd353,
32'sd1935, 32'sd1764, 32'sd148, 32'sd1588, 32'sd1639, 32'sd720,
32'sd110, 32'sd1440, 32'sd218, 32'sd1824, 32'sd975, 32'sd971,
32'sd108, 32'sd1574, 32'sd1042, 32'sd1777, 32'sd870, 32'sd622,
32'sd1846, 32'sd174, 32'sd963, 32'sd651, 32'sd1102, 32'sd136,
32'sd672, 32'sd1553, 32'sd173, 32'sd1437, 32'sd1956, 32'sd593,
32'sd1720, 32'sd762, 32'sd1553, 32'sd801, 32'sd154, 32'sd491,
32'sd1000, 32'sd343, 32'sd627, 32'sd164, 32'sd1298, 32'sd1768,
32'sd1314, 32'sd920, 32'sd669, 32'sd1316, 32'sd1820, 32'sd1315,
32'sd421, 32'sd1970, 32'sd1209, 32'sd1913, 32'sd1771, 32'sd1955,
32'sd1862, 32'sd478, 32'sd956, 32'sd1007, 32'sd647, 32'sd460,
32'sd1881, 32'sd394, 32'sd1598, 32'sd307, 32'sd1333, 32'sd1003,
32'sd1004, 32'sd252, 32'sd1330, 32'sd163, 32'sd1733, 32'sd299,
32'sd1864, 32'sd1024, 32'sd442, 32'sd1991, 32'sd152, 32'sd1406,
32'sd1176, 32'sd1397, 32'sd146, 32'sd1721, 32'sd900, 32'sd1318,
32'sd1700, 32'sd583, 32'sd709, 32'sd1471, 32'sd1448, 32'sd603,
32'sd1476, 32'sd936, 32'sd499, 32'sd1292, 32'sd1810, 32'sd300,
32'sd417, 32'sd1869, 32'sd659, 32'sd974, 32'sd492, 32'sd1516,
32'sd1893, 32'sd1563, 32'sd1182, 32'sd1610, 32'sd446, 32'sd363,
32'sd922, 32'sd1035, 32'sd1274, 32'sd1805, 32'sd1945, 32'sd431,
32'sd1272, 32'sd1940, 32'sd267, 32'sd1181, 32'sd592, 32'sd932,
32'sd1265, 32'sd676, 32'sd316, 32'sd1876, 32'sd1264, 32'sd673,
32'sd1584, 32'sd1573, 32'sd1680, 32'sd343, 32'sd621, 32'sd945,
32'sd1914, 32'sd1434, 32'sd1710, 32'sd581, 32'sd1371, 32'sd1469,
32'sd759, 32'sd1765, 32'sd1177, 32'sd881, 32'sd1455, 32'sd1574,
32'sd682, 32'sd1163, 32'sd1253, 32'sd1251, 32'sd755, 32'sd1423,
32'sd552, 32'sd1889, 32'sd406, 32'sd1693, 32'sd151, 32'sd448,
32'sd1375, 32'sd1408, 32'sd321, 32'sd1841, 32'sd1799, 32'sd1737,
32'sd918, 32'sd1100, 32'sd987, 32'sd807, 32'sd1240, 32'sd718,
32'sd1650, 32'sd1128, 32'sd1201, 32'sd1624, 32'sd776, 32'sd1911,
32'sd476, 32'sd1069, 32'sd942, 32'sd924, 32'sd1845, 32'sd1148,
32'sd846, 32'sd1456, 32'sd1204, 32'sd258, 32'sd321, 32'sd835,
32'sd1789, 32'sd1834, 32'sd1314, 32'sd562, 32'sd1272, 32'sd759,
32'sd1495, 32'sd1289, 32'sd1938, 32'sd1803, 32'sd1937, 32'sd1710,
32'sd845, 32'sd983, 32'sd455, 32'sd1375, 32'sd957, 32'sd1518,
32'sd1951, 32'sd1179, 32'sd1586, 32'sd1012, 32'sd1241, 32'sd1964,
32'sd1881, 32'sd1067, 32'sd1191, 32'sd1141, 32'sd1083, 32'sd1245,
32'sd1878, 32'sd1472, 32'sd1306, 32'sd696, 32'sd143, 32'sd1865,
32'sd1274, 32'sd1647, 32'sd1075, 32'sd1274, 32'sd1189, 32'sd656,
32'sd1944, 32'sd1218, 32'sd931, 32'sd1143, 32'sd1992, 32'sd566,
32'sd1015, 32'sd1773, 32'sd1982, 32'sd456, 32'sd387, 32'sd1091,
32'sd814, 32'sd1209, 32'sd223, 32'sd1240, 32'sd852, 32'sd1178,
32'sd1250, 32'sd1246, 32'sd244, 32'sd693, 32'sd1214, 32'sd198,
32'sd649, 32'sd1949, 32'sd832, 32'sd579, 32'sd1634, 32'sd428,
32'sd748, 32'sd154, 32'sd1363, 32'sd1622, 32'sd1934, 32'sd120,
32'sd243, 32'sd745, 32'sd356, 32'sd712, 32'sd824, 32'sd329,
32'sd988, 32'sd745, 32'sd1321, 32'sd857, 32'sd269, 32'sd1781,
32'sd636, 32'sd1070, 32'sd506, 32'sd1082, 32'sd1981, 32'sd1440,
32'sd647, 32'sd1517, 32'sd437, 32'sd1458, 32'sd708, 32'sd1776,
32'sd1549, 32'sd1658, 32'sd1374, 32'sd204, 32'sd1083, 32'sd939,
32'sd1299, 32'sd1787, 32'sd1282, 32'sd1668, 32'sd1528, 32'sd1287,
32'sd1973, 32'sd996, 32'sd1368, 32'sd1005, 32'sd1388, 32'sd727,
32'sd364, 32'sd1003, 32'sd989, 32'sd1548, 32'sd678, 32'sd1498,
32'sd1761, 32'sd1892, 32'sd161, 32'sd760, 32'sd1969, 32'sd1649,
32'sd1309, 32'sd800, 32'sd529, 32'sd436, 32'sd147, 32'sd1645,
32'sd233, 32'sd773, 32'sd1414, 32'sd1040, 32'sd1798, 32'sd129,
32'sd1294, 32'sd1792, 32'sd1063, 32'sd1485, 32'sd1923, 32'sd1030,
32'sd1556, 32'sd702, 32'sd1012, 32'sd1454, 32'sd116, 32'sd441,
32'sd1904, 32'sd703, 32'sd550, 32'sd235, 32'sd1988, 32'sd1201,
32'sd534, 32'sd1736, 32'sd1823, 32'sd367, 32'sd273, 32'sd1675,
32'sd577, 32'sd796, 32'sd270, 32'sd500, 32'sd1685, 32'sd1691,
32'sd1251, 32'sd521, 32'sd1732, 32'sd1014, 32'sd1291, 32'sd847,
32'sd1811, 32'sd570, 32'sd1587, 32'sd1358, 32'sd1771, 32'sd556,
32'sd1448, 32'sd209, 32'sd1112, 32'sd1978, 32'sd1223, 32'sd1647,
32'sd1643, 32'sd309, 32'sd832, 32'sd389, 32'sd1905, 32'sd1448,
32'sd1266, 32'sd284, 32'sd1610, 32'sd509, 32'sd1119, 32'sd195,
32'sd1799, 32'sd1328, 32'sd1152, 32'sd1029, 32'sd1942, 32'sd737,
32'sd684, 32'sd1319, 32'sd1687, 32'sd1022, 32'sd1863, 32'sd122,
32'sd1761, 32'sd225, 32'sd1763, 32'sd780, 32'sd1906, 32'sd620,
32'sd413, 32'sd1595, 32'sd1666, 32'sd1517, 32'sd938, 32'sd1442,
32'sd1933, 32'sd202, 32'sd101, 32'sd1227, 32'sd1215, 32'sd1891,
32'sd149, 32'sd181, 32'sd1776, 32'sd879, 32'sd608, 32'sd1167,
32'sd1933, 32'sd404, 32'sd1106, 32'sd697, 32'sd561, 32'sd1472,
32'sd1670, 32'sd1395, 32'sd1091, 32'sd371, 32'sd1777, 32'sd199,
32'sd102, 32'sd1532, 32'sd1853, 32'sd1278, 32'sd769, 32'sd1949,
32'sd1230, 32'sd746, 32'sd318, 32'sd1928, 32'sd601, 32'sd1171,
32'sd1766, 32'sd1212, 32'sd956, 32'sd613, 32'sd1294, 32'sd117,
32'sd1048, 32'sd1064, 32'sd952, 32'sd762, 32'sd767, 32'sd614,
32'sd1625, 32'sd1652, 32'sd1156, 32'sd1236, 32'sd1606, 32'sd637,
32'sd572, 32'sd939, 32'sd677, 32'sd726, 32'sd417, 32'sd1299,
32'sd278, 32'sd299, 32'sd278, 32'sd1688, 32'sd596, 32'sd201,
32'sd421, 32'sd742, 32'sd584, 32'sd1878, 32'sd1056, 32'sd1838,
32'sd1617, 32'sd1632, 32'sd1952, 32'sd1246, 32'sd1087, 32'sd1805,
32'sd1106, 32'sd889, 32'sd546, 32'sd1881, 32'sd1561, 32'sd1366,
32'sd483, 32'sd114, 32'sd1207, 32'sd774, 32'sd786, 32'sd1239,
32'sd892, 32'sd505, 32'sd1996, 32'sd596, 32'sd712, 32'sd1808,
32'sd1789, 32'sd1805, 32'sd402, 32'sd1996, 32'sd1941, 32'sd1212,
32'sd1437, 32'sd1732, 32'sd1971, 32'sd1376, 32'sd300, 32'sd1905,
32'sd1477, 32'sd347, 32'sd1770, 32'sd529, 32'sd1154, 32'sd595,
32'sd1077, 32'sd1631, 32'sd1893, 32'sd1357, 32'sd960, 32'sd463,
32'sd973, 32'sd719, 32'sd1289, 32'sd1405, 32'sd530, 32'sd681,
32'sd1256, 32'sd1005, 32'sd1737, 32'sd522, 32'sd1319, 32'sd1450,
32'sd1829, 32'sd1206, 32'sd361, 32'sd953, 32'sd845, 32'sd593,
32'sd1360, 32'sd1249, 32'sd1468, 32'sd1535, 32'sd1959, 32'sd1084,
32'sd1834, 32'sd542, 32'sd473, 32'sd1854, 32'sd1324, 32'sd1961,
32'sd1581, 32'sd744, 32'sd1812, 32'sd1818, 32'sd1474, 32'sd487,
32'sd686, 32'sd1046, 32'sd244, 32'sd116, 32'sd228, 32'sd1670,
32'sd1387, 32'sd237, 32'sd1657, 32'sd1397, 32'sd1149, 32'sd238,
32'sd1521, 32'sd1038, 32'sd1227, 32'sd1880, 32'sd615, 32'sd920,
32'sd1375, 32'sd529, 32'sd934, 32'sd625, 32'sd725, 32'sd181,
32'sd1694, 32'sd1123, 32'sd963, 32'sd619, 32'sd500, 32'sd279,
32'sd902, 32'sd218, 32'sd1004, 32'sd682, 32'sd1495, 32'sd1164,
32'sd454, 32'sd1877, 32'sd560, 32'sd1545, 32'sd1792, 32'sd401,
32'sd332, 32'sd934, 32'sd1215, 32'sd141, 32'sd1199, 32'sd1335,
32'sd1403, 32'sd1393, 32'sd1516, 32'sd1099, 32'sd1216, 32'sd1075,
32'sd814, 32'sd975, 32'sd512, 32'sd1798, 32'sd176, 32'sd151,
32'sd1231, 32'sd1508, 32'sd1810, 32'sd605, 32'sd1358, 32'sd1553,
32'sd633, 32'sd826, 32'sd1004, 32'sd1664, 32'sd735, 32'sd1504,
32'sd218, 32'sd1891, 32'sd1402, 32'sd581, 32'sd105, 32'sd101,
32'sd1686, 32'sd948, 32'sd883, 32'sd578, 32'sd411, 32'sd1100,
32'sd1447, 32'sd1409, 32'sd1592, 32'sd1758, 32'sd118, 32'sd1309,
32'sd1159, 32'sd1983, 32'sd1787, 32'sd1152, 32'sd1129, 32'sd680,
32'sd1067, 32'sd1209, 32'sd666, 32'sd1937, 32'sd1238, 32'sd786,
32'sd1822, 32'sd572, 32'sd263, 32'sd1798, 32'sd1216, 32'sd931,
32'sd1880, 32'sd683, 32'sd1408, 32'sd1736, 32'sd1676, 32'sd419,
32'sd467, 32'sd1915, 32'sd1097, 32'sd795, 32'sd205, 32'sd112,
32'sd128, 32'sd871, 32'sd1028, 32'sd111, 32'sd1712, 32'sd1015,
32'sd353, 32'sd1043, 32'sd513, 32'sd969, 32'sd1419, 32'sd754,
32'sd640, 32'sd1503, 32'sd110, 32'sd806, 32'sd1060, 32'sd579,
32'sd1502, 32'sd1187, 32'sd1624, 32'sd1694, 32'sd821, 32'sd1810,
32'sd683, 32'sd804, 32'sd1356, 32'sd1186, 32'sd1444, 32'sd1324,
32'sd594, 32'sd712, 32'sd1063, 32'sd677, 32'sd614, 32'sd570,
32'sd423, 32'sd1267, 32'sd1177, 32'sd1432, 32'sd1911, 32'sd1554,
32'sd1419, 32'sd731, 32'sd1632, 32'sd1229, 32'sd1343, 32'sd189,
32'sd739, 32'sd952, 32'sd1634, 32'sd128, 32'sd1597, 32'sd1245,
32'sd341, 32'sd1253, 32'sd495, 32'sd1777, 32'sd1731, 32'sd333,
32'sd1408, 32'sd1585, 32'sd145, 32'sd312, 32'sd1735, 32'sd321,
32'sd1071, 32'sd1638, 32'sd221, 32'sd1743, 32'sd158, 32'sd1528,
32'sd1517, 32'sd386, 32'sd927, 32'sd1240, 32'sd1262, 32'sd732,
32'sd1193, 32'sd1508, 32'sd1992, 32'sd189, 32'sd1390, 32'sd1108,
32'sd1337, 32'sd1615, 32'sd797, 32'sd1110, 32'sd1734, 32'sd1880,
32'sd900, 32'sd407, 32'sd1322, 32'sd965, 32'sd406, 32'sd948,
32'sd1278, 32'sd1892, 32'sd1309, 32'sd1417, 32'sd422, 32'sd1300,
32'sd632, 32'sd391, 32'sd1726, 32'sd1270, 32'sd1283, 32'sd1902,
32'sd906, 32'sd1938, 32'sd1741, 32'sd723, 32'sd889, 32'sd1736,
32'sd333, 32'sd197, 32'sd1242, 32'sd586, 32'sd1437, 32'sd583,
32'sd586, 32'sd1058, 32'sd256, 32'sd1793, 32'sd1920, 32'sd1709,
32'sd1422, 32'sd176, 32'sd1076, 32'sd577, 32'sd1037, 32'sd888,
32'sd1046, 32'sd448, 32'sd1340, 32'sd1315, 32'sd1791, 32'sd870,
32'sd1354, 32'sd1892, 32'sd967, 32'sd1001, 32'sd1931, 32'sd842,
32'sd1420, 32'sd615, 32'sd1238, 32'sd1046, 32'sd1291, 32'sd1013,
32'sd314, 32'sd1473, 32'sd1577, 32'sd1951, 32'sd776, 32'sd1445,
32'sd1563, 32'sd105, 32'sd332, 32'sd1271, 32'sd1479, 32'sd1182,
32'sd570, 32'sd1111, 32'sd706, 32'sd154, 32'sd1328, 32'sd1916,
32'sd804, 32'sd1001, 32'sd1056, 32'sd308, 32'sd1914, 32'sd1020,
32'sd1648, 32'sd1992, 32'sd1473, 32'sd1954, 32'sd481, 32'sd300,
32'sd1176, 32'sd1955, 32'sd1900, 32'sd890, 32'sd1701, 32'sd646,
32'sd690, 32'sd1633, 32'sd712, 32'sd1908, 32'sd507, 32'sd1347,
32'sd1600, 32'sd866, 32'sd246, 32'sd1313, 32'sd1489, 32'sd1204,
32'sd1636, 32'sd1416, 32'sd374, 32'sd1011, 32'sd393, 32'sd1144,
32'sd1261, 32'sd903, 32'sd1453, 32'sd816, 32'sd1352, 32'sd180,
32'sd1676, 32'sd867, 32'sd583, 32'sd166, 32'sd1133, 32'sd1510,
32'sd603, 32'sd921, 32'sd543, 32'sd1555, 32'sd952, 32'sd1529,
32'sd1897, 32'sd636, 32'sd407, 32'sd574, 32'sd1560, 32'sd316,
32'sd766, 32'sd1067, 32'sd655, 32'sd1995, 32'sd691, 32'sd402,
32'sd1985, 32'sd340, 32'sd1575, 32'sd115, 32'sd727, 32'sd481,
32'sd955, 32'sd1353, 32'sd831, 32'sd237, 32'sd1408, 32'sd490,
32'sd606, 32'sd655, 32'sd1262, 32'sd1608, 32'sd166, 32'sd257,
32'sd801, 32'sd477, 32'sd226, 32'sd753, 32'sd1151, 32'sd1164,
32'sd688, 32'sd1151, 32'sd1089, 32'sd786, 32'sd1296, 32'sd1254,
32'sd1322, 32'sd847, 32'sd1227, 32'sd365, 32'sd811, 32'sd544,
32'sd1839, 32'sd423, 32'sd1368, 32'sd1394, 32'sd1990, 32'sd1754,
32'sd1622, 32'sd1984, 32'sd543, 32'sd580, 32'sd1606, 32'sd474,
32'sd1399, 32'sd223, 32'sd416, 32'sd1220, 32'sd1167, 32'sd875,
32'sd136, 32'sd576, 32'sd1335, 32'sd656, 32'sd243, 32'sd674,
32'sd951, 32'sd1929, 32'sd1803, 32'sd922, 32'sd1795, 32'sd1993,
32'sd1616, 32'sd1408, 32'sd392, 32'sd1091, 32'sd196, 32'sd1004,
32'sd1321, 32'sd914, 32'sd521, 32'sd1406, 32'sd172, 32'sd680,
32'sd1184, 32'sd1786, 32'sd282, 32'sd152, 32'sd1873, 32'sd808,
32'sd490, 32'sd1306, 32'sd1412, 32'sd1512, 32'sd380, 32'sd768,
32'sd293, 32'sd764, 32'sd1234, 32'sd1740, 32'sd994, 32'sd1399,
32'sd1660, 32'sd904, 32'sd1968, 32'sd1700, 32'sd924, 32'sd486,
32'sd1810, 32'sd1802, 32'sd1155, 32'sd846, 32'sd1480, 32'sd497,
32'sd1890, 32'sd1643, 32'sd1340, 32'sd1435, 32'sd257, 32'sd1560,
32'sd1484, 32'sd1856, 32'sd411, 32'sd908, 32'sd1541, 32'sd358,
32'sd987, 32'sd555, 32'sd802, 32'sd1507, 32'sd1884, 32'sd468,
32'sd814, 32'sd1922, 32'sd1870, 32'sd1267, 32'sd1605, 32'sd410,
32'sd1252, 32'sd1292, 32'sd890, 32'sd263, 32'sd918, 32'sd511,
32'sd1529, 32'sd647, 32'sd1669, 32'sd1906, 32'sd181, 32'sd591,
32'sd1438, 32'sd192, 32'sd564, 32'sd1202, 32'sd1898, 32'sd894,
32'sd1181, 32'sd1759, 32'sd119, 32'sd230, 32'sd1429, 32'sd1907,
32'sd1672, 32'sd829, 32'sd590, 32'sd1201, 32'sd812, 32'sd962,
32'sd1399, 32'sd1751, 32'sd1987, 32'sd717, 32'sd1912, 32'sd593,
32'sd480, 32'sd693, 32'sd1709, 32'sd168, 32'sd1403, 32'sd942,
32'sd1625, 32'sd1185, 32'sd620, 32'sd1116, 32'sd1909, 32'sd1805,
32'sd1523, 32'sd1414, 32'sd504, 32'sd488, 32'sd1775, 32'sd329,
32'sd1639, 32'sd449, 32'sd600, 32'sd1825, 32'sd1187, 32'sd1629,
32'sd877, 32'sd508, 32'sd1902, 32'sd997, 32'sd249, 32'sd1083,
32'sd1238, 32'sd1630, 32'sd137, 32'sd171, 32'sd1040, 32'sd1453,
32'sd1443, 32'sd1964, 32'sd1718, 32'sd813, 32'sd856, 32'sd206,
32'sd525, 32'sd1612, 32'sd1844, 32'sd1893, 32'sd526, 32'sd687,
32'sd1202, 32'sd1667, 32'sd553, 32'sd397, 32'sd624, 32'sd415,
32'sd1892, 32'sd392, 32'sd271, 32'sd406, 32'sd1391, 32'sd691,
32'sd626, 32'sd919, 32'sd775, 32'sd1340, 32'sd1024, 32'sd804,
32'sd709, 32'sd685, 32'sd264, 32'sd1823, 32'sd968, 32'sd1395,
32'sd1514, 32'sd1155, 32'sd1972, 32'sd705, 32'sd1036, 32'sd1275,
32'sd1155, 32'sd1392, 32'sd161, 32'sd661, 32'sd888, 32'sd386,
32'sd735, 32'sd959, 32'sd1983, 32'sd1659, 32'sd1821, 32'sd108,
32'sd1601, 32'sd903, 32'sd1326, 32'sd1376, 32'sd609, 32'sd301,
32'sd657, 32'sd232, 32'sd975, 32'sd1758, 32'sd124, 32'sd113,
32'sd369, 32'sd342, 32'sd1120, 32'sd1802, 32'sd1780, 32'sd140,
32'sd453, 32'sd656, 32'sd725, 32'sd1653, 32'sd1370, 32'sd764,
32'sd317, 32'sd1334, 32'sd380, 32'sd949, 32'sd1033, 32'sd909,
32'sd1577, 32'sd567, 32'sd1035, 32'sd1300, 32'sd217, 32'sd1264,
32'sd282, 32'sd1870, 32'sd749, 32'sd538, 32'sd914, 32'sd171,
32'sd1399, 32'sd1121, 32'sd1126, 32'sd1536, 32'sd1898, 32'sd1679,
32'sd512, 32'sd798, 32'sd1724, 32'sd1521, 32'sd1010, 32'sd1551,
32'sd1391, 32'sd470, 32'sd633, 32'sd1171, 32'sd594, 32'sd1205,
32'sd1755, 32'sd1809, 32'sd472, 32'sd572, 32'sd1944, 32'sd339,
32'sd160, 32'sd1474, 32'sd1919, 32'sd607, 32'sd1275, 32'sd839,
32'sd1839, 32'sd1099, 32'sd500, 32'sd1107, 32'sd1201, 32'sd1556,
32'sd1841, 32'sd495, 32'sd1332, 32'sd2000, 32'sd341, 32'sd1946,
32'sd1184, 32'sd1401, 32'sd271, 32'sd1063, 32'sd815, 32'sd1867,
32'sd1892, 32'sd1790, 32'sd935, 32'sd1697, 32'sd1547, 32'sd1413,
32'sd189, 32'sd1080, 32'sd1580, 32'sd187, 32'sd1087, 32'sd753,
32'sd909, 32'sd106, 32'sd1903, 32'sd1034, 32'sd1243, 32'sd1048,
32'sd719, 32'sd746, 32'sd1807, 32'sd1346, 32'sd257, 32'sd1050,
32'sd1536, 32'sd942, 32'sd1762, 32'sd1720, 32'sd1481, 32'sd1115,
32'sd143, 32'sd711, 32'sd1866, 32'sd472, 32'sd327, 32'sd363,
32'sd532, 32'sd119, 32'sd1891, 32'sd274, 32'sd1231, 32'sd1781,
32'sd664, 32'sd1385, 32'sd668, 32'sd1955, 32'sd1112, 32'sd894,
32'sd166, 32'sd1427, 32'sd1070, 32'sd1928, 32'sd515, 32'sd1539,
32'sd1113, 32'sd725, 32'sd1029, 32'sd1659, 32'sd1006, 32'sd291,
32'sd1786, 32'sd1360, 32'sd768, 32'sd1820, 32'sd107, 32'sd802,
32'sd787, 32'sd1729, 32'sd598, 32'sd722, 32'sd1019, 32'sd1546,
32'sd1432, 32'sd720, 32'sd265, 32'sd167, 32'sd355, 32'sd1871,
32'sd1789, 32'sd587, 32'sd1560, 32'sd1493, 32'sd1014, 32'sd956,
32'sd1094, 32'sd1610, 32'sd1381, 32'sd786, 32'sd535, 32'sd536,
32'sd1654, 32'sd828, 32'sd958, 32'sd1173, 32'sd769, 32'sd1248,
32'sd1544, 32'sd1139, 32'sd1834, 32'sd228, 32'sd976, 32'sd267,
32'sd753, 32'sd411, 32'sd170, 32'sd1197, 32'sd307, 32'sd1890,
32'sd1420, 32'sd900, 32'sd1369, 32'sd903, 32'sd1939, 32'sd1904,
32'sd1088, 32'sd936, 32'sd1475, 32'sd1363, 32'sd584, 32'sd1283,
32'sd1461, 32'sd817, 32'sd1052, 32'sd1489, 32'sd460, 32'sd338,
32'sd1396, 32'sd749, 32'sd1127, 32'sd730, 32'sd1469, 32'sd557,
32'sd1869, 32'sd222, 32'sd1130, 32'sd1928, 32'sd131, 32'sd1205,
32'sd1821, 32'sd604, 32'sd381, 32'sd1532, 32'sd1803, 32'sd1895,
32'sd875, 32'sd1578, 32'sd213, 32'sd674, 32'sd1536, 32'sd633,
32'sd615, 32'sd181, 32'sd1563, 32'sd1257, 32'sd1846, 32'sd121,
32'sd1260, 32'sd1633, 32'sd1342, 32'sd1479, 32'sd1818, 32'sd1703,
32'sd767, 32'sd846, 32'sd167, 32'sd1615, 32'sd1263, 32'sd1237,
32'sd1564, 32'sd640, 32'sd902, 32'sd1951, 32'sd218, 32'sd572,
32'sd620, 32'sd1043, 32'sd1962, 32'sd276, 32'sd1775, 32'sd783,
32'sd481, 32'sd227, 32'sd1485, 32'sd554, 32'sd1672, 32'sd1681,
32'sd1005, 32'sd972, 32'sd411, 32'sd1905, 32'sd919, 32'sd953,
32'sd1125, 32'sd537, 32'sd408, 32'sd670, 32'sd744, 32'sd1330,
32'sd1017, 32'sd1418, 32'sd1553, 32'sd353, 32'sd110, 32'sd417,
32'sd1291, 32'sd1193, 32'sd1153, 32'sd1584, 32'sd1512, 32'sd688,
32'sd657, 32'sd577, 32'sd502, 32'sd1853, 32'sd1712, 32'sd1879,
32'sd889, 32'sd1779, 32'sd1834, 32'sd583, 32'sd1379, 32'sd907,
32'sd268, 32'sd1241, 32'sd807, 32'sd843, 32'sd991, 32'sd1671,
32'sd818, 32'sd800, 32'sd1037, 32'sd1551, 32'sd570, 32'sd122,
32'sd560, 32'sd1298, 32'sd794, 32'sd1686, 32'sd643, 32'sd776,
32'sd635, 32'sd1339, 32'sd1417, 32'sd1651, 32'sd1829, 32'sd965,
32'sd1342, 32'sd242, 32'sd255, 32'sd316, 32'sd1438, 32'sd1243,
32'sd770, 32'sd1467, 32'sd425, 32'sd743, 32'sd838, 32'sd1495,
32'sd163, 32'sd1310, 32'sd355, 32'sd908, 32'sd1908, 32'sd397,
32'sd1193, 32'sd1979, 32'sd694, 32'sd138, 32'sd374, 32'sd955,
32'sd519, 32'sd1171, 32'sd376, 32'sd695, 32'sd1036, 32'sd1977,
32'sd1163, 32'sd1900, 32'sd1843, 32'sd858, 32'sd832, 32'sd1213,
32'sd1395, 32'sd966, 32'sd544, 32'sd356, 32'sd812, 32'sd367,
32'sd781, 32'sd1764, 32'sd842, 32'sd1000, 32'sd1392, 32'sd1011,
32'sd963, 32'sd1292, 32'sd601, 32'sd1963, 32'sd1647, 32'sd1520,
32'sd1718, 32'sd874, 32'sd207, 32'sd1283, 32'sd1566, 32'sd1861,
32'sd192, 32'sd947, 32'sd313, 32'sd870, 32'sd1602, 32'sd1254,
32'sd662, 32'sd1869, 32'sd1368, 32'sd215, 32'sd758, 32'sd1602,
32'sd489, 32'sd863, 32'sd1152, 32'sd912, 32'sd1425, 32'sd1142,
32'sd155, 32'sd716, 32'sd1645, 32'sd1951, 32'sd813, 32'sd108,
32'sd268, 32'sd957, 32'sd666, 32'sd283, 32'sd293, 32'sd1316,
32'sd1335, 32'sd112, 32'sd1152, 32'sd1311, 32'sd912, 32'sd1324,
32'sd1660, 32'sd783, 32'sd975, 32'sd1180, 32'sd1327, 32'sd169,
32'sd1107, 32'sd1441, 32'sd578, 32'sd535, 32'sd148, 32'sd1552,
32'sd1496, 32'sd1433, 32'sd1341, 32'sd1575, 32'sd582, 32'sd694,
32'sd405, 32'sd391, 32'sd1578, 32'sd1937, 32'sd1927, 32'sd897,
32'sd777, 32'sd1348, 32'sd150, 32'sd1799, 32'sd409, 32'sd1527,
32'sd366, 32'sd729, 32'sd1143, 32'sd931, 32'sd515, 32'sd230,
32'sd569, 32'sd1516, 32'sd740, 32'sd1958, 32'sd220, 32'sd1952,
32'sd918, 32'sd942, 32'sd1663, 32'sd503, 32'sd1294, 32'sd966,
32'sd324, 32'sd284, 32'sd1014, 32'sd579, 32'sd665, 32'sd968,
32'sd1588, 32'sd1093, 32'sd1494, 32'sd1272, 32'sd1662, 32'sd377,
32'sd1416, 32'sd105, 32'sd1932, 32'sd367, 32'sd222, 32'sd978,
32'sd781, 32'sd493, 32'sd1968, 32'sd855, 32'sd1192, 32'sd778,
32'sd1362, 32'sd1638, 32'sd103, 32'sd1148, 32'sd1480, 32'sd757,
32'sd955, 32'sd669, 32'sd632, 32'sd581, 32'sd208, 32'sd347,
32'sd1229, 32'sd1481, 32'sd1372, 32'sd693, 32'sd500, 32'sd1199,
32'sd1952, 32'sd1082, 32'sd1451, 32'sd915, 32'sd900, 32'sd717,
32'sd405, 32'sd1119, 32'sd1139, 32'sd1772, 32'sd1004, 32'sd800,
32'sd1540, 32'sd1084, 32'sd553, 32'sd1420, 32'sd359, 32'sd785,
32'sd1363, 32'sd832, 32'sd1662, 32'sd1906, 32'sd448, 32'sd1455,
32'sd567, 32'sd294, 32'sd628, 32'sd1394, 32'sd1492, 32'sd418,
32'sd697, 32'sd276, 32'sd1513, 32'sd1779, 32'sd1980, 32'sd1730,
32'sd1164, 32'sd1160, 32'sd625, 32'sd684, 32'sd955, 32'sd474,
32'sd140, 32'sd768, 32'sd963, 32'sd674, 32'sd634, 32'sd1739,
32'sd1791, 32'sd1442, 32'sd1736, 32'sd1978, 32'sd1592, 32'sd1849,
32'sd1636, 32'sd161, 32'sd578, 32'sd995, 32'sd1685, 32'sd1021,
32'sd1483, 32'sd1748, 32'sd1903, 32'sd599, 32'sd1118, 32'sd714,
32'sd1760, 32'sd1211, 32'sd1552, 32'sd1446, 32'sd801, 32'sd887,
32'sd500, 32'sd967, 32'sd1208, 32'sd360, 32'sd1552, 32'sd844,
32'sd1115, 32'sd931, 32'sd1519, 32'sd1279, 32'sd286, 32'sd665,
32'sd816, 32'sd1552, 32'sd207, 32'sd907, 32'sd1744, 32'sd1040,
32'sd382, 32'sd101, 32'sd547, 32'sd984, 32'sd1186, 32'sd1986,
32'sd1696, 32'sd1433, 32'sd261, 32'sd1456, 32'sd596, 32'sd1358,
32'sd1516, 32'sd1280, 32'sd1768, 32'sd500, 32'sd1873, 32'sd1230,
32'sd170, 32'sd688, 32'sd386, 32'sd1630, 32'sd146, 32'sd1067,
32'sd1210, 32'sd347, 32'sd1977, 32'sd755, 32'sd348, 32'sd1471,
32'sd482, 32'sd1603, 32'sd1555, 32'sd1775, 32'sd328, 32'sd1660,
32'sd1853, 32'sd1322, 32'sd114, 32'sd1198, 32'sd1243, 32'sd1251,
32'sd356, 32'sd1585, 32'sd1331, 32'sd620, 32'sd1306, 32'sd1727,
32'sd540, 32'sd1837, 32'sd586, 32'sd1643, 32'sd1368, 32'sd1502,
32'sd853, 32'sd429, 32'sd994, 32'sd273, 32'sd1139, 32'sd646,
32'sd1560, 32'sd584, 32'sd1524, 32'sd1476, 32'sd361, 32'sd523,
32'sd916, 32'sd1850, 32'sd1885, 32'sd1700, 32'sd200, 32'sd844,
32'sd902, 32'sd312, 32'sd1505, 32'sd847, 32'sd1811, 32'sd820,
32'sd1576, 32'sd1189, 32'sd1516, 32'sd498, 32'sd1110, 32'sd242,
32'sd1344, 32'sd543, 32'sd905, 32'sd904, 32'sd233, 32'sd878,
32'sd426, 32'sd1377, 32'sd218, 32'sd1325, 32'sd646, 32'sd1286,
32'sd479, 32'sd1954, 32'sd195, 32'sd1376, 32'sd1821, 32'sd1366,
32'sd307, 32'sd697, 32'sd481, 32'sd755, 32'sd521, 32'sd923,
32'sd211, 32'sd436, 32'sd1912, 32'sd1334, 32'sd1156, 32'sd907,
32'sd1136, 32'sd1236, 32'sd1648, 32'sd1807, 32'sd1964, 32'sd1814,
32'sd685, 32'sd340, 32'sd1015, 32'sd485, 32'sd106, 32'sd863,
32'sd165, 32'sd251, 32'sd1164, 32'sd289, 32'sd1799, 32'sd1102,
32'sd1518, 32'sd464, 32'sd880, 32'sd671, 32'sd598, 32'sd117,
32'sd1676, 32'sd874, 32'sd329, 32'sd471, 32'sd1421, 32'sd322,
32'sd1552, 32'sd968, 32'sd910, 32'sd1177, 32'sd374, 32'sd555,
32'sd1030, 32'sd710, 32'sd804, 32'sd1213, 32'sd1366, 32'sd1776,
32'sd814, 32'sd1104, 32'sd383, 32'sd987, 32'sd1960, 32'sd1327,
32'sd1724, 32'sd1263, 32'sd1890, 32'sd664, 32'sd1649, 32'sd924,
32'sd930, 32'sd1661, 32'sd1607, 32'sd1221, 32'sd1133, 32'sd1506,
32'sd1191, 32'sd1902, 32'sd1395, 32'sd1786, 32'sd268, 32'sd410,
32'sd316, 32'sd1813, 32'sd1811, 32'sd1354, 32'sd181, 32'sd1976,
32'sd601, 32'sd1289, 32'sd345, 32'sd581, 32'sd375, 32'sd1033,
32'sd1777, 32'sd1554, 32'sd1971, 32'sd1592, 32'sd469, 32'sd192,
32'sd139, 32'sd1554, 32'sd1729, 32'sd162, 32'sd1410, 32'sd1833,
32'sd1221, 32'sd577, 32'sd1635, 32'sd867, 32'sd1005, 32'sd137,
32'sd409, 32'sd1680, 32'sd918, 32'sd1363, 32'sd581, 32'sd1469,
32'sd922, 32'sd1902, 32'sd683, 32'sd1296, 32'sd1018, 32'sd1016,
32'sd1788, 32'sd1224, 32'sd1100, 32'sd1831, 32'sd1966, 32'sd394,
32'sd824, 32'sd1185, 32'sd1814, 32'sd571, 32'sd1851, 32'sd1917,
32'sd836, 32'sd1908, 32'sd1152, 32'sd553, 32'sd758, 32'sd687,
32'sd402, 32'sd950, 32'sd162, 32'sd753, 32'sd1384, 32'sd602,
32'sd1473, 32'sd1737, 32'sd1637, 32'sd631, 32'sd363, 32'sd471,
32'sd1493, 32'sd297, 32'sd1203, 32'sd1820, 32'sd958, 32'sd1061,
32'sd124, 32'sd1197, 32'sd281, 32'sd1699, 32'sd1714, 32'sd854,
32'sd566, 32'sd517, 32'sd245, 32'sd1184, 32'sd1613, 32'sd1270,
32'sd1315, 32'sd1026, 32'sd1195, 32'sd219, 32'sd1544, 32'sd1330,
32'sd433, 32'sd1647, 32'sd261, 32'sd306, 32'sd556, 32'sd1606,
32'sd929, 32'sd995, 32'sd1195, 32'sd1403, 32'sd1270, 32'sd373,
32'sd1261, 32'sd248, 32'sd1852, 32'sd1389, 32'sd1891, 32'sd1855,
32'sd918, 32'sd1109, 32'sd1598, 32'sd656, 32'sd546, 32'sd692,
32'sd400, 32'sd392, 32'sd132, 32'sd1137, 32'sd795, 32'sd1878,
32'sd662, 32'sd1643, 32'sd820, 32'sd832, 32'sd1526, 32'sd1959,
32'sd105, 32'sd1475, 32'sd150, 32'sd1579, 32'sd1217, 32'sd1389,
32'sd779, 32'sd349, 32'sd1275, 32'sd892, 32'sd599, 32'sd190,
32'sd1610, 32'sd1261, 32'sd1259, 32'sd855, 32'sd673, 32'sd1053,
32'sd1782, 32'sd1675, 32'sd1315, 32'sd484, 32'sd927, 32'sd522,
32'sd1779, 32'sd1932, 32'sd333, 32'sd1331, 32'sd1757, 32'sd1475,
32'sd461, 32'sd1808, 32'sd595, 32'sd1418, 32'sd1915, 32'sd1942,
32'sd489, 32'sd1605, 32'sd801, 32'sd633, 32'sd975, 32'sd518,
32'sd800, 32'sd1709, 32'sd1429, 32'sd1470, 32'sd816, 32'sd132,
32'sd171, 32'sd1296, 32'sd1041, 32'sd630, 32'sd704, 32'sd575,
32'sd966, 32'sd1892, 32'sd751, 32'sd910, 32'sd1105, 32'sd633,
32'sd428, 32'sd593, 32'sd1276, 32'sd1312, 32'sd899, 32'sd1405,
32'sd643, 32'sd1099, 32'sd1035, 32'sd308, 32'sd707, 32'sd1748,
32'sd1255, 32'sd926, 32'sd657, 32'sd1520, 32'sd503, 32'sd1451,
32'sd794, 32'sd1368, 32'sd1860, 32'sd816, 32'sd1838, 32'sd1349,
32'sd207, 32'sd1320, 32'sd1653, 32'sd134, 32'sd1116, 32'sd862,
32'sd353, 32'sd912, 32'sd1664, 32'sd1762, 32'sd431, 32'sd1864,
32'sd1472, 32'sd590, 32'sd726, 32'sd1618, 32'sd919, 32'sd1248,
32'sd194, 32'sd1737, 32'sd905, 32'sd1390, 32'sd1156, 32'sd1485,
32'sd1641, 32'sd251, 32'sd402, 32'sd1887, 32'sd1857, 32'sd307,
32'sd334, 32'sd1041, 32'sd906, 32'sd400, 32'sd1374, 32'sd191,
32'sd1693, 32'sd1660, 32'sd154, 32'sd584, 32'sd1070, 32'sd1903,
32'sd927, 32'sd125, 32'sd1891, 32'sd207, 32'sd1761, 32'sd1591,
32'sd777, 32'sd1744, 32'sd156, 32'sd192, 32'sd1942, 32'sd842,
32'sd1098, 32'sd1526, 32'sd636, 32'sd1099, 32'sd1623, 32'sd1577,
32'sd659, 32'sd1293, 32'sd165, 32'sd1766, 32'sd701, 32'sd1256,
32'sd799, 32'sd568, 32'sd1640, 32'sd150, 32'sd770, 32'sd331,
32'sd202, 32'sd254, 32'sd1150, 32'sd1906, 32'sd140, 32'sd878,
32'sd278, 32'sd1636, 32'sd1881, 32'sd919, 32'sd1167, 32'sd1955,
32'sd1510, 32'sd712, 32'sd934, 32'sd1229, 32'sd1415, 32'sd852,
32'sd793, 32'sd1313, 32'sd1160, 32'sd389, 32'sd464, 32'sd1323,
32'sd620, 32'sd333, 32'sd968, 32'sd810, 32'sd240, 32'sd1866,
32'sd1953, 32'sd757, 32'sd863, 32'sd1580, 32'sd1517, 32'sd1765,
32'sd1826, 32'sd1610, 32'sd792, 32'sd1856, 32'sd1397, 32'sd1199,
32'sd1286, 32'sd377, 32'sd1209, 32'sd1854, 32'sd1955, 32'sd280,
32'sd1874, 32'sd1030, 32'sd1281, 32'sd1234, 32'sd1257, 32'sd425,
32'sd639, 32'sd709, 32'sd808, 32'sd619, 32'sd1660, 32'sd1044,
32'sd1573, 32'sd1039, 32'sd1773, 32'sd1312, 32'sd1070, 32'sd1334,
32'sd233, 32'sd1719, 32'sd1094, 32'sd1167, 32'sd1213, 32'sd1839,
32'sd437, 32'sd729, 32'sd1188, 32'sd1379, 32'sd707, 32'sd1951,
32'sd1358, 32'sd215, 32'sd753, 32'sd179, 32'sd1202, 32'sd644,
32'sd738, 32'sd1823, 32'sd199, 32'sd632, 32'sd504, 32'sd242,
32'sd166, 32'sd1253, 32'sd1547, 32'sd264, 32'sd1338, 32'sd1856,
32'sd1482, 32'sd1538, 32'sd398, 32'sd1730, 32'sd423, 32'sd228,
32'sd195, 32'sd1524, 32'sd630, 32'sd1640, 32'sd1636, 32'sd798,
32'sd1412, 32'sd1591, 32'sd327, 32'sd108, 32'sd1695, 32'sd961,
32'sd1776, 32'sd1002, 32'sd1776, 32'sd463, 32'sd758, 32'sd1995,
32'sd469, 32'sd1903, 32'sd1995, 32'sd921, 32'sd1850, 32'sd992,
32'sd441, 32'sd1789, 32'sd490, 32'sd1362, 32'sd1054, 32'sd1862,
32'sd1204, 32'sd632, 32'sd411, 32'sd1413, 32'sd526, 32'sd1077,
32'sd1515, 32'sd792, 32'sd1671, 32'sd1436, 32'sd1700, 32'sd957,
32'sd445, 32'sd1329, 32'sd546, 32'sd1497, 32'sd1423, 32'sd1794,
32'sd1208, 32'sd1946, 32'sd388, 32'sd1268, 32'sd274, 32'sd1088,
32'sd1089, 32'sd1404, 32'sd1077, 32'sd448, 32'sd1798, 32'sd791,
32'sd1455, 32'sd1251, 32'sd702, 32'sd1914, 32'sd1060, 32'sd1841,
32'sd1930, 32'sd1724, 32'sd679, 32'sd337, 32'sd1175, 32'sd1087,
32'sd1017, 32'sd1036, 32'sd691, 32'sd1681, 32'sd862, 32'sd869,
32'sd374, 32'sd243, 32'sd328, 32'sd1664, 32'sd1697, 32'sd452,
32'sd1525, 32'sd1120, 32'sd570, 32'sd1331, 32'sd1313, 32'sd258,
32'sd1278, 32'sd1532, 32'sd1920, 32'sd1617, 32'sd1423, 32'sd1806,
32'sd1119, 32'sd1744, 32'sd1516, 32'sd650, 32'sd392, 32'sd1274,
32'sd137, 32'sd1076, 32'sd1354, 32'sd727, 32'sd668, 32'sd586,
32'sd489, 32'sd1064, 32'sd666, 32'sd587, 32'sd714, 32'sd275,
32'sd1314, 32'sd320, 32'sd1650, 32'sd1389, 32'sd871, 32'sd444,
32'sd393, 32'sd129, 32'sd186, 32'sd321, 32'sd1828, 32'sd1157,
32'sd1848, 32'sd1908, 32'sd1955, 32'sd1346, 32'sd1561, 32'sd1711,
32'sd549, 32'sd1689, 32'sd1763, 32'sd1908, 32'sd1715, 32'sd1560,
32'sd1800, 32'sd477, 32'sd1553, 32'sd1895, 32'sd612, 32'sd728,
32'sd1118, 32'sd931, 32'sd931, 32'sd1903, 32'sd572, 32'sd1403,
32'sd276, 32'sd568, 32'sd1118, 32'sd112, 32'sd1370, 32'sd1265,
32'sd1483, 32'sd340, 32'sd1101, 32'sd1966, 32'sd741, 32'sd1638,
32'sd789, 32'sd1499, 32'sd320, 32'sd145, 32'sd276, 32'sd790,
32'sd430, 32'sd1485, 32'sd543, 32'sd1991, 32'sd143, 32'sd1893,
32'sd1494, 32'sd1954, 32'sd262, 32'sd1160, 32'sd410, 32'sd956,
32'sd1754, 32'sd659, 32'sd758, 32'sd378, 32'sd341, 32'sd1801,
32'sd1916, 32'sd1721, 32'sd1218, 32'sd1205, 32'sd1451, 32'sd934,
32'sd381, 32'sd929, 32'sd1271, 32'sd609, 32'sd1470, 32'sd1690,
32'sd1374, 32'sd550, 32'sd1616, 32'sd929, 32'sd1263, 32'sd1374,
32'sd1500, 32'sd1946, 32'sd541, 32'sd535, 32'sd920, 32'sd1846,
32'sd1838, 32'sd968, 32'sd744, 32'sd1861, 32'sd1907, 32'sd924,
32'sd271, 32'sd1596, 32'sd113, 32'sd1629, 32'sd1819, 32'sd1762,
32'sd1161, 32'sd1047, 32'sd1340, 32'sd836, 32'sd1647, 32'sd1187,
32'sd1196, 32'sd1638, 32'sd1542, 32'sd167, 32'sd128, 32'sd1253,
32'sd499, 32'sd1243, 32'sd1481, 32'sd1947, 32'sd1954, 32'sd1851,
32'sd1626, 32'sd1164, 32'sd1327, 32'sd942, 32'sd1023, 32'sd1927
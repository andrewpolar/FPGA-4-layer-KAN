32'sd1128711, 32'sd786731,
32'sd507842, 32'sd510350,
32'sd858079, 32'sd1174114,
32'sd599110, 32'sd563914,
32'sd732518, 32'sd617970,
32'sd778122, 32'sd885450,
32'sd759075, 32'sd643785,
32'sd847802, 32'sd668559,
32'sd612115, 32'sd783834,
32'sd967588, 32'sd860088,
32'sd525597, 32'sd1125088,
32'sd1167246, 32'sd509733,
32'sd647029, 32'sd801035,
32'sd858613, 32'sd983999,
32'sd841815, 32'sd1154688,
32'sd1174309, 32'sd477543,
32'sd1067995, 32'sd1200838,
32'sd1039374, 32'sd1128600,
32'sd1146863, 32'sd1042500,
32'sd692088, 32'sd1035171,
32'sd1016393, 32'sd1002968,
32'sd976651, 32'sd748269,
32'sd920111, 32'sd697179,
32'sd709321, 32'sd507875,
32'sd915195, 32'sd529053,
32'sd1130344, 32'sd865901,
32'sd1178849, 32'sd1028142,
32'sd726183, 32'sd589734,
32'sd1175508, 32'sd1130679,
32'sd1039756, 32'sd452190,
32'sd692044, 32'sd743572,
32'sd738458, 32'sd702351,
32'sd676504, 32'sd985301,
32'sd484285, 32'sd1193261,
32'sd640468, 32'sd993068,
32'sd1187299, 32'sd601333,
32'sd739712, 32'sd914997,
32'sd972329, 32'sd856689,
32'sd925364, 32'sd557223,
32'sd759649, 32'sd878404,
32'sd691486, 32'sd739370,
32'sd549567, 32'sd1208543,
32'sd1055977, 32'sd646276,
32'sd1006149, 32'sd848449,
32'sd831394, 32'sd709081,
32'sd496039, 32'sd846420,
32'sd863571, 32'sd830664,
32'sd628319, 32'sd1026134,
32'sd506978, 32'sd405403,
32'sd959976, 32'sd590051,
32'sd876951, 32'sd465775,
32'sd829474, 32'sd886140,
32'sd554196, 32'sd1009181,
32'sd831345, 32'sd501252,
32'sd537923, 32'sd910900,
32'sd977087, 32'sd802120,
32'sd945268, 32'sd948455,
32'sd773860, 32'sd987595,
32'sd1006178, 32'sd584974,
32'sd1125916, 32'sd834064,
32'sd733861, 32'sd618198,
32'sd769188, 32'sd800102,
32'sd575220, 32'sd1033196,
32'sd421924, 32'sd761875,
32'sd428767, 32'sd801919,
32'sd718022, 32'sd804403,
32'sd938332, 32'sd1139635,
32'sd972732, 32'sd433998,
32'sd664819, 32'sd1116935,
32'sd1165633, 32'sd1168514,
32'sd1127207, 32'sd907542,
32'sd679600, 32'sd1072753,
32'sd1053191, 32'sd1201577,
32'sd1045977, 32'sd503723,
32'sd920910, 32'sd459199,
32'sd600538, 32'sd1064442,
32'sd666917, 32'sd976591,
32'sd839859, 32'sd582060,
32'sd759959, 32'sd530129,
32'sd805543, 32'sd505036,
32'sd626759, 32'sd1174973,
32'sd713005, 32'sd1111607,
32'sd922604, 32'sd1107359,
32'sd863023, 32'sd931499,
32'sd533705, 32'sd1037882,
32'sd1124220, 32'sd639708,
32'sd823450, 32'sd812578,
32'sd662445, 32'sd462513,
32'sd1118824, 32'sd1145223,
32'sd804623, 32'sd1185853,
32'sd924000, 32'sd947719,
32'sd982063, 32'sd456768,
32'sd763381, 32'sd770661,
32'sd711355, 32'sd687476,
32'sd675428, 32'sd601509,
32'sd573287, 32'sd814034,
32'sd845962, 32'sd764241,
32'sd1091673, 32'sd739871,
32'sd1064143, 32'sd1059888,
32'sd523589, 32'sd507168,
32'sd819255, 32'sd729089,
32'sd1115485, 32'sd477337,
32'sd506778, 32'sd796749,
32'sd424751, 32'sd969660,
32'sd1034103, 32'sd418973,
32'sd872846, 32'sd841421,
32'sd1158452, 32'sd1142553,
32'sd983646, 32'sd817161,
32'sd640144, 32'sd1159140,
32'sd837190, 32'sd652329,
32'sd632901, 32'sd469588,
32'sd932594, 32'sd1007668,
32'sd949469, 32'sd575240,
32'sd621784, 32'sd468534,
32'sd697521, 32'sd909634,
32'sd911915, 32'sd511078,
32'sd633377, 32'sd1061243,
32'sd852545, 32'sd1009485,
32'sd913193, 32'sd874769,
32'sd975774, 32'sd941809,
32'sd470123, 32'sd1057772,
32'sd1177250, 32'sd751844,
32'sd485178, 32'sd1043446,
32'sd916809, 32'sd910916,
32'sd843806, 32'sd758032,
32'sd524187, 32'sd1204516,
32'sd887943, 32'sd690844,
32'sd1020373, 32'sd482072,
32'sd706616, 32'sd965139,
32'sd824152, 32'sd626141,
32'sd751741, 32'sd880290,
32'sd469581, 32'sd663578,
32'sd753042, 32'sd410702,
32'sd833590, 32'sd1204295,
32'sd592547, 32'sd1195895,
32'sd897430, 32'sd934515,
32'sd1119448, 32'sd527260,
32'sd668595, 32'sd571772,
32'sd772838, 32'sd584130,
32'sd1190078, 32'sd958516,
32'sd1105319, 32'sd647878,
32'sd1138633, 32'sd1161001,
32'sd708829, 32'sd923258,
32'sd631916, 32'sd1078113,
32'sd480951, 32'sd729829,
32'sd1126823, 32'sd1123439,
32'sd427482, 32'sd943148,
32'sd675279, 32'sd766620,
32'sd507900, 32'sd785110,
32'sd1043217, 32'sd1017887,
32'sd704572, 32'sd552105,
32'sd1059410, 32'sd1087767,
32'sd731400, 32'sd558652,
32'sd731520, 32'sd791286,
32'sd1036210, 32'sd421357,
32'sd1183058, 32'sd661200,
32'sd1189280, 32'sd1144017,
32'sd1072424, 32'sd1004531,
32'sd477773, 32'sd989492,
32'sd647981, 32'sd760941,
32'sd1074163, 32'sd469811,
32'sd597109, 32'sd441407,
32'sd1099826, 32'sd433720,
32'sd636885, 32'sd985669,
32'sd1136608, 32'sd995770,
32'sd556967, 32'sd725941,
32'sd1133815, 32'sd466684,
32'sd663472, 32'sd1124151,
32'sd494090, 32'sd550533,
32'sd667649, 32'sd690661,
32'sd1114501, 32'sd683345,
32'sd1022596, 32'sd1062525,
32'sd1154073, 32'sd439438,
32'sd537192, 32'sd1044069,
32'sd1118918, 32'sd509764,
32'sd552707, 32'sd687197,
32'sd786964, 32'sd756249,
32'sd642288, 32'sd753644,
32'sd618519, 32'sd510860,
32'sd852800, 32'sd568583,
32'sd617306, 32'sd1133914,
32'sd763486, 32'sd791141,
32'sd594317, 32'sd501729,
32'sd492048, 32'sd982325,
32'sd689622, 32'sd1042374,
32'sd673019, 32'sd666696,
32'sd624530, 32'sd677186,
32'sd1025098, 32'sd615234,
32'sd728846, 32'sd848546,
32'sd579978, 32'sd1066009,
32'sd491325, 32'sd840574,
32'sd1119464, 32'sd487470,
32'sd1104479, 32'sd700219,
32'sd1065145, 32'sd1159627,
32'sd735255, 32'sd744519,
32'sd872979, 32'sd582101,
32'sd1000661, 32'sd1164888,
32'sd678696, 32'sd795166,
32'sd1123914, 32'sd801562,
32'sd817079, 32'sd880082,
32'sd932714, 32'sd411531,
32'sd436893, 32'sd499686,
32'sd589052, 32'sd1104411,
32'sd530204, 32'sd1096477,
32'sd1188145, 32'sd1174128,
32'sd846066, 32'sd972564,
32'sd1058989, 32'sd495823,
32'sd1014920, 32'sd688423,
32'sd837050, 32'sd1062543,
32'sd1046662, 32'sd1180564,
32'sd548414, 32'sd520539,
32'sd848725, 32'sd772422,
32'sd594408, 32'sd542142,
32'sd1094626, 32'sd692108,
32'sd1080848, 32'sd687111,
32'sd933945, 32'sd759694,
32'sd614097, 32'sd779977,
32'sd1178531, 32'sd1118262,
32'sd457727, 32'sd1209811,
32'sd924212, 32'sd1010000,
32'sd701452, 32'sd444720,
32'sd428061, 32'sd682945,
32'sd973510, 32'sd526950,
32'sd640609, 32'sd901655,
32'sd1164825, 32'sd758178,
32'sd612439, 32'sd615797,
32'sd656467, 32'sd730516,
32'sd535044, 32'sd623983,
32'sd817695, 32'sd921651,
32'sd683608, 32'sd791770,
32'sd963311, 32'sd1023069,
32'sd561808, 32'sd718837,
32'sd852804, 32'sd1104328,
32'sd499499, 32'sd441217,
32'sd685311, 32'sd689863,
32'sd726808, 32'sd422811,
32'sd801137, 32'sd798328,
32'sd598372, 32'sd449161,
32'sd520483, 32'sd728704,
32'sd886469, 32'sd884689,
32'sd684465, 32'sd687467,
32'sd641674, 32'sd605255,
32'sd587015, 32'sd914395,
32'sd463861, 32'sd516602,
32'sd538157, 32'sd910908,
32'sd740265, 32'sd1181556,
32'sd747234, 32'sd887379,
32'sd1019770, 32'sd791341,
32'sd981536, 32'sd1137541,
32'sd675228, 32'sd656858,
32'sd557198, 32'sd1151402,
32'sd615728, 32'sd535320,
32'sd533967, 32'sd1002320,
32'sd878144, 32'sd588904,
32'sd917601, 32'sd1073076,
32'sd526589, 32'sd800716,
32'sd869993, 32'sd1070489,
32'sd822107, 32'sd760804,
32'sd1132025, 32'sd458291,
32'sd1012191, 32'sd870600,
32'sd772539, 32'sd498538,
32'sd979585, 32'sd1132591,
32'sd636274, 32'sd994993,
32'sd1131511, 32'sd904750,
32'sd816594, 32'sd841114,
32'sd543619, 32'sd1073937,
32'sd1152534, 32'sd850988,
32'sd1093384, 32'sd810276,
32'sd425581, 32'sd667243,
32'sd901132, 32'sd1014086,
32'sd1068122, 32'sd1006959,
32'sd821166, 32'sd1111223,
32'sd755685, 32'sd1045710,
32'sd605734, 32'sd1162928,
32'sd1115917, 32'sd833214,
32'sd806914, 32'sd1060113,
32'sd823395, 32'sd546329,
32'sd1033679, 32'sd427345,
32'sd942470, 32'sd536406,
32'sd517211, 32'sd830889,
32'sd512435, 32'sd1195098,
32'sd1070226, 32'sd847527,
32'sd1109590, 32'sd951602,
32'sd1191426, 32'sd426140,
32'sd457861, 32'sd1169908,
32'sd1037904, 32'sd737369,
32'sd979808, 32'sd569514,
32'sd872395, 32'sd974950,
32'sd531938, 32'sd844515,
32'sd706953, 32'sd607046,
32'sd602055, 32'sd1190039,
32'sd793907, 32'sd919868,
32'sd1064327, 32'sd475408,
32'sd643810, 32'sd698745,
32'sd1023988, 32'sd1031041,
32'sd508126, 32'sd775514,
32'sd552413, 32'sd1052437,
32'sd830642, 32'sd458948,
32'sd1111372, 32'sd419024,
32'sd765382, 32'sd1036199,
32'sd691126, 32'sd629680,
32'sd1101524, 32'sd1138806,
32'sd1180253, 32'sd964795,
32'sd695520, 32'sd483906,
32'sd1139700, 32'sd967572,
32'sd573212, 32'sd712409,
32'sd989969, 32'sd716150,
32'sd497058, 32'sd428349,
32'sd1132344, 32'sd637917,
32'sd1148923, 32'sd1168765,
32'sd411945, 32'sd544338,
32'sd544897, 32'sd579658,
32'sd1170373, 32'sd1084634,
32'sd647105, 32'sd1151220,
32'sd746124, 32'sd1162752,
32'sd855313, 32'sd576452,
32'sd1092299, 32'sd934877,
32'sd834752, 32'sd635574
32'sd616217, 32'sd797751, 32'sd994240, 32'sd913779, 32'sd963522, 32'sd828513, 32'sd868514, 32'sd595420, 32'sd519635, 32'sd1189702, 32'sd965239, 32'sd1123674, 32'sd903071, 32'sd1158742,
32'sd942045, 32'sd809807, 32'sd542854, 32'sd919236, 32'sd564453, 32'sd452141, 32'sd921536, 32'sd1198309, 32'sd597739, 32'sd835086, 32'sd1158050, 32'sd787062, 32'sd792937, 32'sd910244,
32'sd976397, 32'sd571238, 32'sd1196582, 32'sd422420, 32'sd451145, 32'sd770698, 32'sd698125, 32'sd1101428, 32'sd793980, 32'sd757867, 32'sd1035209, 32'sd1103678, 32'sd886646, 32'sd545834,
32'sd1060894, 32'sd631525, 32'sd410508, 32'sd686817, 32'sd581016, 32'sd408347, 32'sd722841, 32'sd628674, 32'sd839534, 32'sd406092, 32'sd1097685, 32'sd920067, 32'sd1188259, 32'sd1140290,
32'sd1037531, 32'sd899746, 32'sd1155914, 32'sd442726, 32'sd868697, 32'sd660045, 32'sd738800, 32'sd558736, 32'sd886429, 32'sd998472, 32'sd867350, 32'sd916297, 32'sd1060619, 32'sd1137362,
32'sd978182, 32'sd975188, 32'sd1044250, 32'sd498898, 32'sd509786, 32'sd965529, 32'sd607282, 32'sd880440, 32'sd1143183, 32'sd451694, 32'sd1105467, 32'sd624591, 32'sd652623, 32'sd1183345,
32'sd509498, 32'sd492837, 32'sd554196, 32'sd1030743, 32'sd925118, 32'sd663094, 32'sd487945, 32'sd612230, 32'sd742437, 32'sd450353, 32'sd744380, 32'sd429324, 32'sd635669, 32'sd641738,
32'sd1071126, 32'sd431974, 32'sd1039180, 32'sd888339, 32'sd1113032, 32'sd464389, 32'sd910236, 32'sd1173868, 32'sd1205241, 32'sd644197, 32'sd789984, 32'sd1147425, 32'sd578547, 32'sd1026694,
32'sd502279, 32'sd1113279, 32'sd487839, 32'sd702550, 32'sd705245, 32'sd884475, 32'sd1132495, 32'sd671632, 32'sd851053, 32'sd817814, 32'sd853215, 32'sd956228, 32'sd1202705, 32'sd1100914,
32'sd1037952, 32'sd580106, 32'sd1157878, 32'sd472462, 32'sd1158570, 32'sd830474, 32'sd518962, 32'sd798057, 32'sd462818, 32'sd529643, 32'sd1192157, 32'sd744814, 32'sd664770, 32'sd1027430,
32'sd1154500, 32'sd680763, 32'sd982588, 32'sd946629, 32'sd671266, 32'sd668510, 32'sd1194027, 32'sd935842, 32'sd583982, 32'sd749508, 32'sd421007, 32'sd989953, 32'sd912768, 32'sd863080,
32'sd598773, 32'sd593258, 32'sd1138829, 32'sd462874, 32'sd715809, 32'sd528566, 32'sd651730, 32'sd859445, 32'sd526919, 32'sd1110102, 32'sd757953, 32'sd554122, 32'sd1063908, 32'sd1041355,
32'sd1042197, 32'sd764053, 32'sd1097499, 32'sd1127012, 32'sd935237, 32'sd1171417, 32'sd661693, 32'sd1188391, 32'sd497186, 32'sd507707, 32'sd989171, 32'sd673338, 32'sd1086927, 32'sd537915,
32'sd1026217, 32'sd768872, 32'sd773848, 32'sd597966, 32'sd834481, 32'sd438026, 32'sd714499, 32'sd1121867, 32'sd497571, 32'sd639695, 32'sd893617, 32'sd658862, 32'sd642043, 32'sd726199,
32'sd726552, 32'sd776834, 32'sd434442, 32'sd619849, 32'sd1079968, 32'sd982089, 32'sd623817, 32'sd759349, 32'sd792672, 32'sd960861, 32'sd1205073, 32'sd859328, 32'sd875713, 32'sd1041703,
32'sd1181880, 32'sd936915, 32'sd866555, 32'sd591690, 32'sd480621, 32'sd778755, 32'sd527773, 32'sd618585, 32'sd1193080, 32'sd935485, 32'sd990784, 32'sd1104286, 32'sd863944, 32'sd655249,
32'sd763973, 32'sd960331, 32'sd627889, 32'sd630509, 32'sd1177386, 32'sd1100845, 32'sd1056251, 32'sd1196762, 32'sd1207788, 32'sd822832, 32'sd414275, 32'sd1179391, 32'sd631008, 32'sd421180,
32'sd544735, 32'sd1026299, 32'sd603208, 32'sd602954, 32'sd491106, 32'sd1003953, 32'sd765129, 32'sd418611, 32'sd1114210, 32'sd1155832, 32'sd685696, 32'sd1001975, 32'sd1185103, 32'sd996071,
32'sd928285, 32'sd1001918, 32'sd410813, 32'sd910838, 32'sd1155332, 32'sd794532, 32'sd595310, 32'sd995735, 32'sd602066, 32'sd659968, 32'sd564939, 32'sd522711, 32'sd637812, 32'sd1124197,
32'sd504806, 32'sd571690, 32'sd1013151, 32'sd829873, 32'sd1089462, 32'sd811577, 32'sd1135653, 32'sd815287, 32'sd666710, 32'sd597669, 32'sd1129588, 32'sd1100140, 32'sd1015375, 32'sd476994,
32'sd1114689, 32'sd536302, 32'sd1090778, 32'sd436124, 32'sd705459, 32'sd451756, 32'sd690559, 32'sd834448, 32'sd428805, 32'sd1073229, 32'sd407420, 32'sd485274, 32'sd489511, 32'sd727333,
32'sd717833, 32'sd419668, 32'sd754332, 32'sd776254, 32'sd708339, 32'sd523331, 32'sd527835, 32'sd692124, 32'sd1116045, 32'sd689473, 32'sd1150989, 32'sd954719, 32'sd716944, 32'sd419652,
32'sd1156730, 32'sd867849, 32'sd1032072, 32'sd1077166, 32'sd951261, 32'sd567555, 32'sd595540, 32'sd1071506, 32'sd1182148, 32'sd498390, 32'sd1109318, 32'sd472802, 32'sd476758, 32'sd811769,
32'sd1205618, 32'sd777173, 32'sd565915, 32'sd777110, 32'sd876012, 32'sd892957, 32'sd1046565, 32'sd880045, 32'sd621211, 32'sd978952, 32'sd434937, 32'sd930683, 32'sd769519, 32'sd1182293,
32'sd1161974, 32'sd798845, 32'sd524845, 32'sd1004469, 32'sd546799, 32'sd606702, 32'sd1180322, 32'sd1091705, 32'sd562947, 32'sd598279, 32'sd546646, 32'sd531934, 32'sd818008, 32'sd624896,
32'sd1111423, 32'sd429906, 32'sd517154, 32'sd925747, 32'sd813749, 32'sd764879, 32'sd577264, 32'sd501596, 32'sd477274, 32'sd743863, 32'sd994433, 32'sd1122244, 32'sd596811, 32'sd788310,
32'sd732628, 32'sd529866, 32'sd1183809, 32'sd1048776, 32'sd488113, 32'sd1182671, 32'sd998157, 32'sd1002055, 32'sd629754, 32'sd570677, 32'sd1158558, 32'sd659047, 32'sd994131, 32'sd904233,
32'sd980123, 32'sd1144548, 32'sd698851, 32'sd917064, 32'sd1171679, 32'sd979918, 32'sd848953, 32'sd985184, 32'sd741485, 32'sd1198001, 32'sd543754, 32'sd1164105, 32'sd528221, 32'sd1119654,
32'sd428843, 32'sd686980, 32'sd564403, 32'sd1113208, 32'sd612624, 32'sd530684, 32'sd679042, 32'sd605674, 32'sd817458, 32'sd934442, 32'sd435721, 32'sd1205320, 32'sd938157, 32'sd713554,
32'sd1032387, 32'sd828563, 32'sd1152458, 32'sd924063, 32'sd935540, 32'sd962539, 32'sd815725, 32'sd781314, 32'sd1113282, 32'sd551870, 32'sd1122727, 32'sd1075544, 32'sd675901, 32'sd1176901,
32'sd1092993, 32'sd414176, 32'sd656474, 32'sd549145, 32'sd675215, 32'sd893427, 32'sd1167457, 32'sd616627, 32'sd1110600, 32'sd1117576, 32'sd434090, 32'sd961618, 32'sd427572, 32'sd947737,
32'sd847165, 32'sd1059034, 32'sd482561, 32'sd667492, 32'sd1016028, 32'sd1178091, 32'sd1144763, 32'sd647612, 32'sd1096039, 32'sd726892, 32'sd681601, 32'sd679859, 32'sd442985, 32'sd677368,
32'sd1121328, 32'sd671717, 32'sd918391, 32'sd689885, 32'sd978194, 32'sd600068, 32'sd450263, 32'sd1068527, 32'sd743395, 32'sd885579, 32'sd852652, 32'sd724038, 32'sd1168055, 32'sd1094270,
32'sd705086, 32'sd668721, 32'sd970973, 32'sd1064753, 32'sd1098588, 32'sd548781, 32'sd440361, 32'sd1002702, 32'sd520190, 32'sd804735, 32'sd1017248, 32'sd736387, 32'sd685662, 32'sd1025168,
32'sd780808, 32'sd1161284, 32'sd442338, 32'sd536831, 32'sd854292, 32'sd513402, 32'sd988668, 32'sd817607, 32'sd829957, 32'sd990626, 32'sd460250, 32'sd578490, 32'sd803991, 32'sd1002025,
32'sd453819, 32'sd1048585, 32'sd528795, 32'sd638697, 32'sd613591, 32'sd597395, 32'sd709537, 32'sd847925, 32'sd503891, 32'sd492875, 32'sd900758, 32'sd468286, 32'sd589307, 32'sd591429,
32'sd436563, 32'sd758416, 32'sd1187154, 32'sd867955, 32'sd851944, 32'sd1184682, 32'sd945560, 32'sd593486, 32'sd1155338, 32'sd413952, 32'sd578963, 32'sd606255, 32'sd962370, 32'sd872009,
32'sd933578, 32'sd514160, 32'sd738072, 32'sd1007965, 32'sd640218, 32'sd915131, 32'sd766557, 32'sd513731, 32'sd417697, 32'sd525346, 32'sd459255, 32'sd858433, 32'sd537732, 32'sd434961,
32'sd533883, 32'sd534224, 32'sd1005783, 32'sd896649, 32'sd1018635, 32'sd786612, 32'sd671095, 32'sd891704, 32'sd827920, 32'sd611203, 32'sd1192500, 32'sd1016087, 32'sd639738, 32'sd701265,
32'sd1039386, 32'sd1024760, 32'sd1120328, 32'sd1085951, 32'sd560774, 32'sd756389, 32'sd428486, 32'sd612955, 32'sd784809, 32'sd892276, 32'sd994653, 32'sd958786, 32'sd453174, 32'sd482462,
32'sd404614, 32'sd430338, 32'sd1078859, 32'sd983206, 32'sd1094132, 32'sd428358, 32'sd714963, 32'sd695559, 32'sd499376, 32'sd607286, 32'sd1010808, 32'sd1087090, 32'sd986398, 32'sd824364,
32'sd947496, 32'sd1171511, 32'sd685219, 32'sd1023118, 32'sd507782, 32'sd1092212, 32'sd947157, 32'sd703527, 32'sd471399, 32'sd653535, 32'sd463975, 32'sd783633, 32'sd927811, 32'sd475961,
32'sd558867, 32'sd1001998, 32'sd958477, 32'sd1005290, 32'sd986141, 32'sd665415, 32'sd1019819, 32'sd676117, 32'sd1208141, 32'sd923749, 32'sd417732, 32'sd1104532, 32'sd874278, 32'sd445852,
32'sd436671, 32'sd1025666, 32'sd889921, 32'sd537114, 32'sd984103, 32'sd458085, 32'sd961033, 32'sd484941, 32'sd873693, 32'sd779733, 32'sd662420, 32'sd690890, 32'sd457787, 32'sd462519,
32'sd1047324, 32'sd780204, 32'sd410362, 32'sd741945, 32'sd642712, 32'sd889711, 32'sd611968, 32'sd1081974, 32'sd897456, 32'sd439082, 32'sd1079888, 32'sd1075769, 32'sd737635, 32'sd446554,
32'sd829687, 32'sd584830, 32'sd490710, 32'sd885111, 32'sd948253, 32'sd997817, 32'sd972213, 32'sd639567, 32'sd526596, 32'sd953230, 32'sd573199, 32'sd1059821, 32'sd687866, 32'sd896270,
32'sd1096428, 32'sd1106639, 32'sd976709, 32'sd434948, 32'sd1022205, 32'sd819916, 32'sd540668, 32'sd407203, 32'sd505310, 32'sd510196, 32'sd675203, 32'sd724555, 32'sd1186746, 32'sd850658,
32'sd674843, 32'sd524580, 32'sd1068009, 32'sd515566, 32'sd1167056, 32'sd467990, 32'sd786001, 32'sd791890, 32'sd584127, 32'sd863946, 32'sd732809, 32'sd944495, 32'sd809804, 32'sd1029957,
32'sd843844, 32'sd1125138, 32'sd471705, 32'sd592671, 32'sd610666, 32'sd812798, 32'sd779648, 32'sd1125853, 32'sd663553, 32'sd1014656, 32'sd964180, 32'sd555664, 32'sd1019950, 32'sd1128798,
32'sd1082985, 32'sd713469, 32'sd475945, 32'sd471914, 32'sd462116, 32'sd763196, 32'sd680202, 32'sd1018511, 32'sd1019638, 32'sd819836, 32'sd1025653, 32'sd805852, 32'sd1124686, 32'sd812401,
32'sd935679, 32'sd569063, 32'sd538014, 32'sd680878, 32'sd802758, 32'sd1062824, 32'sd406228, 32'sd618185, 32'sd538003, 32'sd700373, 32'sd756030, 32'sd1018109, 32'sd607206, 32'sd1065628,
32'sd875014, 32'sd1068450, 32'sd1002045, 32'sd593051, 32'sd1164484, 32'sd497717, 32'sd574895, 32'sd444511, 32'sd625350, 32'sd778795, 32'sd844196, 32'sd1015779, 32'sd443397, 32'sd507936,
32'sd1033263, 32'sd948148, 32'sd441136, 32'sd1198075, 32'sd1196222, 32'sd573308, 32'sd464092, 32'sd890147, 32'sd854143, 32'sd1064023, 32'sd913250, 32'sd1158140, 32'sd875409, 32'sd1059650,
32'sd897902, 32'sd589121, 32'sd781983, 32'sd888612, 32'sd924908, 32'sd696925, 32'sd1073731, 32'sd857447, 32'sd668849, 32'sd1197911, 32'sd418060, 32'sd1120490, 32'sd893758, 32'sd858450,
32'sd808008, 32'sd611250, 32'sd777180, 32'sd973363, 32'sd1174842, 32'sd579473, 32'sd758029, 32'sd789133, 32'sd950816, 32'sd826987, 32'sd1159375, 32'sd723724, 32'sd627815, 32'sd1207483,
32'sd585258, 32'sd570048, 32'sd821906, 32'sd600455, 32'sd807478, 32'sd1072418, 32'sd789380, 32'sd1162228, 32'sd439459, 32'sd889459, 32'sd516420, 32'sd702149, 32'sd580863, 32'sd939454,
32'sd544299, 32'sd1154908, 32'sd503006, 32'sd696664, 32'sd749873, 32'sd1155447, 32'sd795234, 32'sd966360, 32'sd1007330, 32'sd521747, 32'sd777753, 32'sd621398, 32'sd1117082, 32'sd779151,
32'sd842812, 32'sd688637, 32'sd779007, 32'sd776596, 32'sd482152, 32'sd1071398, 32'sd758479, 32'sd1188611, 32'sd822462, 32'sd1075760, 32'sd971124, 32'sd1003655, 32'sd451310, 32'sd1034594,
32'sd978508, 32'sd1030803, 32'sd1103004, 32'sd983097, 32'sd1082786, 32'sd772933, 32'sd743149, 32'sd587000, 32'sd616576, 32'sd544253, 32'sd1161236, 32'sd1059586, 32'sd1155646, 32'sd702329,
32'sd908976, 32'sd915550, 32'sd640556, 32'sd463627, 32'sd1060796, 32'sd818225, 32'sd1028454, 32'sd581820, 32'sd753345, 32'sd589679, 32'sd538593, 32'sd445570, 32'sd783573, 32'sd551738,
32'sd1085087, 32'sd773688, 32'sd1081160, 32'sd459376, 32'sd904444, 32'sd999971, 32'sd467119, 32'sd1176849, 32'sd1122658, 32'sd1148251, 32'sd522779, 32'sd974849, 32'sd923758, 32'sd1148854,
32'sd435147, 32'sd1131224, 32'sd1164442, 32'sd1195616, 32'sd1167945, 32'sd745768, 32'sd1012733, 32'sd832835, 32'sd939268, 32'sd969225, 32'sd769268, 32'sd600501, 32'sd616562, 32'sd699551,
32'sd496568, 32'sd698899, 32'sd1083596, 32'sd1016436, 32'sd451537, 32'sd501596, 32'sd730263, 32'sd1130207, 32'sd573736, 32'sd664933, 32'sd746521, 32'sd543966, 32'sd1034913, 32'sd712071,
32'sd1202997, 32'sd437258, 32'sd406051, 32'sd461511, 32'sd670271, 32'sd799869, 32'sd646856, 32'sd677310, 32'sd830595, 32'sd588244, 32'sd895103, 32'sd854992, 32'sd1121895, 32'sd704116,
32'sd1127378, 32'sd433241, 32'sd538950, 32'sd1079834, 32'sd567864, 32'sd1120810, 32'sd550801, 32'sd525060, 32'sd824319, 32'sd899544, 32'sd678214, 32'sd725721, 32'sd900589, 32'sd978751,
32'sd848222, 32'sd981787, 32'sd582392, 32'sd788019, 32'sd1193960, 32'sd555517, 32'sd1169464, 32'sd518389, 32'sd659417, 32'sd749521, 32'sd666075, 32'sd1088531, 32'sd502335, 32'sd929892,
32'sd426045, 32'sd440961, 32'sd648608, 32'sd480007, 32'sd537603, 32'sd1195769, 32'sd663741, 32'sd442554, 32'sd829793, 32'sd1172344, 32'sd1171129, 32'sd890036, 32'sd1089384, 32'sd562518,
32'sd753566, 32'sd468990, 32'sd721107, 32'sd580119, 32'sd534918, 32'sd1126359, 32'sd785040, 32'sd889343, 32'sd579058, 32'sd553798, 32'sd753198, 32'sd1168058, 32'sd594490, 32'sd593117,
32'sd756987, 32'sd492074, 32'sd471738, 32'sd1145618, 32'sd828019, 32'sd1153879, 32'sd648270, 32'sd416948, 32'sd705561, 32'sd955473, 32'sd1084925, 32'sd840472, 32'sd614035, 32'sd1200766,
32'sd1186996, 32'sd794494, 32'sd980732, 32'sd448454, 32'sd1179360, 32'sd894536, 32'sd770205, 32'sd1192807, 32'sd1070989, 32'sd934646, 32'sd703984, 32'sd924762, 32'sd519636, 32'sd1148430,
32'sd1156382, 32'sd428082, 32'sd1027135, 32'sd759509, 32'sd879495, 32'sd434599, 32'sd880809, 32'sd817215, 32'sd941773, 32'sd746929, 32'sd541434, 32'sd414125, 32'sd963207, 32'sd850781,
32'sd576234, 32'sd806020, 32'sd1047058, 32'sd748011, 32'sd684958, 32'sd728854, 32'sd789234, 32'sd935477, 32'sd469791, 32'sd480338, 32'sd1207710, 32'sd1158180, 32'sd849243, 32'sd501221,
32'sd1139265, 32'sd630770, 32'sd861216, 32'sd1105629, 32'sd1129612, 32'sd498979, 32'sd1172126, 32'sd1067842, 32'sd560211, 32'sd1151057, 32'sd620681, 32'sd1034454, 32'sd512231, 32'sd1013377,
32'sd797893, 32'sd1020094, 32'sd1173228, 32'sd695567, 32'sd476064, 32'sd814886, 32'sd1102286, 32'sd466584, 32'sd846641, 32'sd856378, 32'sd868192, 32'sd760928, 32'sd881484, 32'sd745978,
32'sd900220, 32'sd710438, 32'sd485846, 32'sd1068963, 32'sd793391, 32'sd816870, 32'sd951368, 32'sd477689, 32'sd544491, 32'sd601339, 32'sd408530, 32'sd457221, 32'sd520323, 32'sd1055515,
32'sd879805, 32'sd682204, 32'sd489571, 32'sd1182097, 32'sd1013223, 32'sd505260, 32'sd988227, 32'sd535362, 32'sd560693, 32'sd850044, 32'sd688183, 32'sd951039, 32'sd489756, 32'sd1113314,
32'sd761705, 32'sd1053386, 32'sd943527, 32'sd553079, 32'sd860468, 32'sd1125753, 32'sd792317, 32'sd976089, 32'sd974132, 32'sd506038, 32'sd480397, 32'sd1035445, 32'sd612072, 32'sd623020,
32'sd721447, 32'sd913180, 32'sd1126344, 32'sd505909, 32'sd489744, 32'sd451049, 32'sd938781, 32'sd410125, 32'sd1151937, 32'sd1146991, 32'sd576524, 32'sd747777, 32'sd1120750, 32'sd1031714,
32'sd1169807, 32'sd1195831, 32'sd752860, 32'sd1159458, 32'sd456094, 32'sd744746, 32'sd818696, 32'sd1158830, 32'sd917040, 32'sd1062016, 32'sd1128113, 32'sd478513, 32'sd693124, 32'sd1064033,
32'sd541975, 32'sd620611, 32'sd801120, 32'sd1180941, 32'sd873966, 32'sd1107667, 32'sd1089778, 32'sd707184, 32'sd590469, 32'sd771282, 32'sd754874, 32'sd564828, 32'sd447007, 32'sd1112203,
32'sd570971, 32'sd458798, 32'sd627857, 32'sd1086223, 32'sd1126113, 32'sd1069449, 32'sd779294, 32'sd547897, 32'sd610423, 32'sd1178612, 32'sd976000, 32'sd815512, 32'sd405271, 32'sd426173,
32'sd967643, 32'sd770499, 32'sd603294, 32'sd816950, 32'sd1038281, 32'sd953818, 32'sd1085753, 32'sd730476, 32'sd807852, 32'sd1184217, 32'sd801060, 32'sd918919, 32'sd626967, 32'sd598035,
32'sd428389, 32'sd455425, 32'sd587437, 32'sd714538, 32'sd1171892, 32'sd895113, 32'sd629559, 32'sd680533, 32'sd536036, 32'sd894222, 32'sd603597, 32'sd987446, 32'sd936212, 32'sd960802,
32'sd869533, 32'sd683662, 32'sd633868, 32'sd723524, 32'sd456302, 32'sd1145188, 32'sd798510, 32'sd450227, 32'sd738611, 32'sd795855, 32'sd935476, 32'sd811219, 32'sd1050557, 32'sd579184,
32'sd628279, 32'sd699164, 32'sd404402, 32'sd679649, 32'sd692717, 32'sd898273, 32'sd1084601, 32'sd1023882, 32'sd1017899, 32'sd780680, 32'sd1094371, 32'sd653826, 32'sd567146, 32'sd1033993,
32'sd1052773, 32'sd1103344, 32'sd505213, 32'sd1210049, 32'sd470389, 32'sd936970, 32'sd953246, 32'sd1072687, 32'sd1134472, 32'sd1135194, 32'sd805252, 32'sd683393, 32'sd553754, 32'sd1125268,
32'sd778383, 32'sd995563, 32'sd642571, 32'sd980809, 32'sd476441, 32'sd498619, 32'sd935380, 32'sd922488, 32'sd996015, 32'sd512375, 32'sd514900, 32'sd1196419, 32'sd1071093, 32'sd685941,
32'sd1203794, 32'sd605382, 32'sd563372, 32'sd621439, 32'sd1132970, 32'sd1153190, 32'sd785315, 32'sd1085159, 32'sd1081392, 32'sd594968, 32'sd661483, 32'sd1125965, 32'sd824530, 32'sd571227,
32'sd527710, 32'sd442253, 32'sd814426, 32'sd816741, 32'sd632598, 32'sd822314, 32'sd510480, 32'sd520619, 32'sd765921, 32'sd707318, 32'sd998541, 32'sd518078, 32'sd797915, 32'sd1077768,
32'sd632259, 32'sd705760, 32'sd403975, 32'sd794800, 32'sd1200136, 32'sd910484, 32'sd430370, 32'sd732252, 32'sd632038, 32'sd795645, 32'sd867437, 32'sd1031654, 32'sd678957, 32'sd783515,
32'sd918319, 32'sd1204397, 32'sd1145511, 32'sd975228, 32'sd852116, 32'sd1041057, 32'sd750926, 32'sd638793, 32'sd619239, 32'sd647350, 32'sd624738, 32'sd454458, 32'sd671512, 32'sd1031000,
32'sd579942, 32'sd498801, 32'sd877884, 32'sd872806, 32'sd625250, 32'sd481383, 32'sd499240, 32'sd1002828, 32'sd406634, 32'sd864521, 32'sd888159, 32'sd1165626, 32'sd679840, 32'sd910106,
32'sd900688, 32'sd517549, 32'sd457241, 32'sd752157, 32'sd563293, 32'sd1134083, 32'sd489633, 32'sd1000062, 32'sd710452, 32'sd749834, 32'sd735176, 32'sd430549, 32'sd913225, 32'sd1169678,
32'sd1178635, 32'sd889473, 32'sd900877, 32'sd563153, 32'sd648362, 32'sd1113604, 32'sd797361, 32'sd860426, 32'sd506998, 32'sd476706, 32'sd651764, 32'sd737634, 32'sd805038, 32'sd704206,
32'sd1017816, 32'sd766230, 32'sd1076047, 32'sd768494, 32'sd585497, 32'sd1058158, 32'sd616144, 32'sd531502, 32'sd1038930, 32'sd1081325, 32'sd1047416, 32'sd1077995, 32'sd540961, 32'sd892715,
32'sd1206066, 32'sd959294, 32'sd855778, 32'sd473975, 32'sd985833, 32'sd540224, 32'sd1066235, 32'sd863801, 32'sd687711, 32'sd598528, 32'sd688476, 32'sd970752, 32'sd434654, 32'sd965620,
32'sd902215, 32'sd417929, 32'sd488238, 32'sd801476, 32'sd1194775, 32'sd747495, 32'sd437815, 32'sd856744, 32'sd977763, 32'sd505001, 32'sd1117280, 32'sd852416, 32'sd1007491, 32'sd512324,
32'sd821281, 32'sd1163560, 32'sd813352, 32'sd905037, 32'sd972382, 32'sd942309, 32'sd824185, 32'sd1088630, 32'sd423195, 32'sd730697, 32'sd624230, 32'sd709388, 32'sd840127, 32'sd648725,
32'sd1144972, 32'sd840270, 32'sd864346, 32'sd720725, 32'sd1193905, 32'sd540538, 32'sd482130, 32'sd430456, 32'sd527149, 32'sd446076, 32'sd961121, 32'sd613612, 32'sd544239, 32'sd774982,
32'sd1051719, 32'sd1191846, 32'sd1134247, 32'sd874741, 32'sd493113, 32'sd1124688, 32'sd1137482, 32'sd629595, 32'sd647849, 32'sd1148700, 32'sd492581, 32'sd821597, 32'sd494513, 32'sd781859,
32'sd823185, 32'sd935538, 32'sd578673, 32'sd739204, 32'sd754956, 32'sd1015727, 32'sd510853, 32'sd1025581, 32'sd1191877, 32'sd1022309, 32'sd824316, 32'sd936188, 32'sd792489, 32'sd884818,
32'sd913386, 32'sd909875, 32'sd1207336, 32'sd1103757, 32'sd1024604, 32'sd1003895, 32'sd864562, 32'sd511163, 32'sd412701, 32'sd827271, 32'sd1033570, 32'sd497028, 32'sd1121878, 32'sd819093,
32'sd1170274, 32'sd1167512, 32'sd1149762, 32'sd1176361, 32'sd951258, 32'sd618860, 32'sd820752, 32'sd631798, 32'sd481446, 32'sd938135, 32'sd497119, 32'sd892997, 32'sd658658, 32'sd635350,
32'sd817680, 32'sd781717, 32'sd810414, 32'sd552991, 32'sd590424, 32'sd909061, 32'sd736369, 32'sd733303, 32'sd1096216, 32'sd852989, 32'sd565248, 32'sd1159558, 32'sd642025, 32'sd944573,
32'sd579190, 32'sd975834, 32'sd582276, 32'sd697097, 32'sd771425, 32'sd954699, 32'sd1007128, 32'sd695039, 32'sd689443, 32'sd1051034, 32'sd801413, 32'sd444716, 32'sd858671, 32'sd1054905,
32'sd939642, 32'sd459800, 32'sd629371, 32'sd508899, 32'sd648080, 32'sd991937, 32'sd1108820, 32'sd947586, 32'sd1105057, 32'sd563744, 32'sd677767, 32'sd740025, 32'sd727519, 32'sd867642,
32'sd1186644, 32'sd1192785, 32'sd599985, 32'sd1033952, 32'sd421694, 32'sd1123755, 32'sd1047709, 32'sd734662, 32'sd910485, 32'sd1134757, 32'sd852575, 32'sd1062067, 32'sd1080117, 32'sd1093296,
32'sd832297, 32'sd735437, 32'sd1011286, 32'sd907508, 32'sd753883, 32'sd1072055, 32'sd415356, 32'sd651269, 32'sd1203553, 32'sd796146, 32'sd1145598, 32'sd1180252, 32'sd672802, 32'sd1205196,
32'sd436060, 32'sd901877, 32'sd627696, 32'sd769968, 32'sd466299, 32'sd982870, 32'sd797206, 32'sd976051, 32'sd766494, 32'sd919859, 32'sd569827, 32'sd787517, 32'sd593318, 32'sd797713,
32'sd1114558, 32'sd788140, 32'sd565370, 32'sd652684, 32'sd1051067, 32'sd555729, 32'sd983181, 32'sd1164131, 32'sd745258, 32'sd1123068, 32'sd732788, 32'sd877909, 32'sd730906, 32'sd841783,
32'sd1039491, 32'sd930842, 32'sd811088, 32'sd1036219, 32'sd931046, 32'sd803268, 32'sd1203664, 32'sd975492, 32'sd849570, 32'sd1163643, 32'sd612597, 32'sd929197, 32'sd1061854, 32'sd944876,
32'sd1171796, 32'sd757919, 32'sd893869, 32'sd605251, 32'sd610510, 32'sd633432, 32'sd616343, 32'sd831961, 32'sd898663, 32'sd527565, 32'sd583305, 32'sd1176441, 32'sd982919, 32'sd580860,
32'sd500462, 32'sd674323, 32'sd968356, 32'sd649117, 32'sd848416, 32'sd1059429, 32'sd743045, 32'sd1200021, 32'sd1067010, 32'sd1093912, 32'sd592493, 32'sd725796, 32'sd478407, 32'sd995419,
32'sd915480, 32'sd571914, 32'sd540688, 32'sd976486, 32'sd457465, 32'sd537479, 32'sd470042, 32'sd1084805, 32'sd791539, 32'sd593482, 32'sd1062606, 32'sd432496, 32'sd671027, 32'sd411740,
32'sd987818, 32'sd639940, 32'sd1174946, 32'sd679618, 32'sd1061877, 32'sd1167176, 32'sd950738, 32'sd446945, 32'sd1142112, 32'sd832133, 32'sd808496, 32'sd646299, 32'sd808650, 32'sd593215,
32'sd726216, 32'sd1088573, 32'sd767336, 32'sd1047244, 32'sd912843, 32'sd560438, 32'sd614449, 32'sd799420, 32'sd594130, 32'sd1094975, 32'sd775930, 32'sd692599, 32'sd405366, 32'sd982846,
32'sd558196, 32'sd931776, 32'sd803774, 32'sd741778, 32'sd1153991, 32'sd768767, 32'sd1039806, 32'sd588651, 32'sd1193044, 32'sd491756, 32'sd420678, 32'sd915436, 32'sd458934, 32'sd626203,
32'sd1044570, 32'sd492075, 32'sd944523, 32'sd555331, 32'sd611155, 32'sd1058530, 32'sd575140, 32'sd518634, 32'sd533814, 32'sd724302, 32'sd1200434, 32'sd1077940, 32'sd820202, 32'sd730526,
32'sd953664, 32'sd1177928, 32'sd983567, 32'sd871585, 32'sd1136840, 32'sd831208, 32'sd945286, 32'sd675335, 32'sd684912, 32'sd495480, 32'sd1180717, 32'sd498108, 32'sd709491, 32'sd905782,
32'sd555596, 32'sd1059880, 32'sd933071, 32'sd871792, 32'sd754541, 32'sd918003, 32'sd411428, 32'sd424583, 32'sd657699, 32'sd657151, 32'sd1143770, 32'sd719534, 32'sd931270, 32'sd1177308,
32'sd1098840, 32'sd687769, 32'sd1028667, 32'sd892046, 32'sd559505, 32'sd780301, 32'sd459463, 32'sd1019926, 32'sd773169, 32'sd523312, 32'sd570057, 32'sd758880, 32'sd712430, 32'sd1090354,
32'sd581012, 32'sd927907, 32'sd741111, 32'sd897223, 32'sd582318, 32'sd645002, 32'sd495310, 32'sd943765, 32'sd544326, 32'sd1109184, 32'sd707857, 32'sd502363, 32'sd858577, 32'sd549803,
32'sd610695, 32'sd466885, 32'sd416692, 32'sd900682, 32'sd643817, 32'sd1055484, 32'sd771801, 32'sd965370, 32'sd991446, 32'sd877646, 32'sd1137321, 32'sd587058, 32'sd416681, 32'sd654995,
32'sd1041537, 32'sd650164, 32'sd682877, 32'sd847931, 32'sd804423, 32'sd439219, 32'sd727575, 32'sd984146, 32'sd647646, 32'sd1054059, 32'sd621626, 32'sd859506, 32'sd747201, 32'sd899682,
32'sd571194, 32'sd426135, 32'sd991073, 32'sd932999, 32'sd787578, 32'sd1025661, 32'sd1077707, 32'sd409567, 32'sd712805, 32'sd567208, 32'sd1089346, 32'sd711855, 32'sd776124, 32'sd534938,
32'sd1049077, 32'sd586203, 32'sd439053, 32'sd922856, 32'sd555574, 32'sd911847, 32'sd458326, 32'sd1172790, 32'sd739692, 32'sd1021653, 32'sd808096, 32'sd900727, 32'sd978118, 32'sd511420,
32'sd1139671, 32'sd905269, 32'sd1127632, 32'sd622642, 32'sd783792, 32'sd782841, 32'sd479990, 32'sd979067, 32'sd783484, 32'sd1058760, 32'sd690684, 32'sd1133934, 32'sd1048317, 32'sd567465,
32'sd989216, 32'sd608062, 32'sd647123, 32'sd984014, 32'sd1063478, 32'sd602907, 32'sd508553, 32'sd1155233, 32'sd759874, 32'sd887062, 32'sd665621, 32'sd1137343, 32'sd564439, 32'sd550288,
32'sd1106012, 32'sd1081648, 32'sd1186451, 32'sd651500, 32'sd466912, 32'sd1152716, 32'sd577686, 32'sd787958, 32'sd428329, 32'sd1099676, 32'sd624054, 32'sd775914, 32'sd712147, 32'sd483831,
32'sd557017, 32'sd813530, 32'sd968263, 32'sd726806, 32'sd701875, 32'sd999055, 32'sd880925, 32'sd1127679, 32'sd802153, 32'sd500060, 32'sd801331, 32'sd1161547, 32'sd845062, 32'sd714699,
32'sd887904, 32'sd821496, 32'sd873152, 32'sd1040072, 32'sd796950, 32'sd1175205, 32'sd650374, 32'sd1041114, 32'sd999977, 32'sd577448, 32'sd793592, 32'sd758726, 32'sd513231, 32'sd996015,
32'sd1043852, 32'sd1184155, 32'sd841646, 32'sd1153345, 32'sd513247, 32'sd743954, 32'sd1153582, 32'sd991411, 32'sd621623, 32'sd684841, 32'sd443862, 32'sd410115, 32'sd1172335, 32'sd1207118,
32'sd545938, 32'sd563874, 32'sd653089, 32'sd709824, 32'sd551719, 32'sd1077024, 32'sd514543, 32'sd904898, 32'sd758011, 32'sd883584, 32'sd414071, 32'sd1053732, 32'sd765572, 32'sd1027897,
32'sd676790, 32'sd1060675, 32'sd632329, 32'sd943090, 32'sd622060, 32'sd725947, 32'sd639045, 32'sd969002, 32'sd931388, 32'sd1189761, 32'sd776409, 32'sd954804, 32'sd481999, 32'sd560756,
32'sd446008, 32'sd918437, 32'sd554243, 32'sd531989, 32'sd506481, 32'sd683843, 32'sd857193, 32'sd1017327, 32'sd599709, 32'sd987271, 32'sd989195, 32'sd468839, 32'sd842577, 32'sd695475,
32'sd760442, 32'sd1102926, 32'sd825797, 32'sd681969, 32'sd967548, 32'sd942098, 32'sd446135, 32'sd423463, 32'sd476897, 32'sd712166, 32'sd450551, 32'sd472039, 32'sd1122723, 32'sd1169966,
32'sd714275, 32'sd882939, 32'sd562856, 32'sd1155886, 32'sd889216, 32'sd893743, 32'sd523039, 32'sd749304, 32'sd455368, 32'sd947628, 32'sd741451, 32'sd1116711, 32'sd430402, 32'sd842270,
32'sd776312, 32'sd758309, 32'sd942099, 32'sd1061883, 32'sd1077685, 32'sd1115496, 32'sd415271, 32'sd883584, 32'sd824316, 32'sd610414, 32'sd798393, 32'sd869109, 32'sd478247, 32'sd1046005,
32'sd1003050, 32'sd627810, 32'sd967400, 32'sd453194, 32'sd1123638, 32'sd1173507, 32'sd555119, 32'sd549984, 32'sd436585, 32'sd513685, 32'sd889856, 32'sd634161, 32'sd919964, 32'sd1069405,
32'sd1079225, 32'sd513589, 32'sd621771, 32'sd740453, 32'sd565516, 32'sd992970, 32'sd549721, 32'sd772670, 32'sd763214, 32'sd448194, 32'sd543633, 32'sd710164, 32'sd636849, 32'sd867615,
32'sd1106251, 32'sd996725, 32'sd1110152, 32'sd1125768, 32'sd837629, 32'sd821717, 32'sd449275, 32'sd588380, 32'sd875586, 32'sd1053151, 32'sd1203838, 32'sd513443, 32'sd503370, 32'sd589496,
32'sd486926, 32'sd816560, 32'sd757433, 32'sd1161791, 32'sd448570, 32'sd907124, 32'sd429931, 32'sd1087015, 32'sd1168072, 32'sd675639, 32'sd954394, 32'sd1197375, 32'sd1084859, 32'sd1067520,
32'sd732608, 32'sd603538, 32'sd950386, 32'sd476503, 32'sd796730, 32'sd875085, 32'sd925038, 32'sd861109, 32'sd601427, 32'sd984157, 32'sd1035612, 32'sd1148078, 32'sd939680, 32'sd460669,
32'sd751148, 32'sd710373, 32'sd1085261, 32'sd1125798, 32'sd1140285, 32'sd751234, 32'sd893720, 32'sd992420, 32'sd932990, 32'sd1182891, 32'sd1095401, 32'sd924119, 32'sd1200633, 32'sd917069,
32'sd672586, 32'sd1074866, 32'sd423512, 32'sd1134708, 32'sd803014, 32'sd414070, 32'sd843861, 32'sd1060580, 32'sd1112833, 32'sd735000, 32'sd532747, 32'sd467809, 32'sd422377, 32'sd654185,
32'sd761854, 32'sd885363, 32'sd1171043, 32'sd877094, 32'sd1002790, 32'sd501813, 32'sd859764, 32'sd519202, 32'sd983245, 32'sd1095686, 32'sd1186509, 32'sd882481, 32'sd947445, 32'sd758473,
32'sd660466, 32'sd468854, 32'sd1197004, 32'sd947457, 32'sd871255, 32'sd997172, 32'sd587367, 32'sd773971, 32'sd497137, 32'sd958788, 32'sd583618, 32'sd512463, 32'sd708302, 32'sd824177,
32'sd977025, 32'sd811869, 32'sd1026316, 32'sd589076, 32'sd1033679, 32'sd1066200, 32'sd613898, 32'sd1207764, 32'sd598303, 32'sd856912, 32'sd1065842, 32'sd536584, 32'sd742820, 32'sd691439,
32'sd866985, 32'sd584574, 32'sd525793, 32'sd604719, 32'sd449661, 32'sd923372, 32'sd587996, 32'sd528896, 32'sd564315, 32'sd886146, 32'sd944304, 32'sd517431, 32'sd533509, 32'sd1023827,
32'sd1008812, 32'sd514880, 32'sd910948, 32'sd999530, 32'sd882998, 32'sd427400, 32'sd454258, 32'sd514124, 32'sd961749, 32'sd704162, 32'sd1163676, 32'sd1185618, 32'sd479529, 32'sd582014,
32'sd833136, 32'sd1090310, 32'sd466300, 32'sd521216, 32'sd639742, 32'sd415322, 32'sd580701, 32'sd960001, 32'sd629379, 32'sd422013, 32'sd932515, 32'sd900929, 32'sd851500, 32'sd630962,
32'sd744001, 32'sd982088, 32'sd769877, 32'sd1202133, 32'sd747499, 32'sd1168754, 32'sd1116966, 32'sd936607, 32'sd1026772, 32'sd648218, 32'sd446000, 32'sd1142595, 32'sd966418, 32'sd551715,
32'sd1074608, 32'sd1043413, 32'sd653784, 32'sd1003815, 32'sd595080, 32'sd819896, 32'sd1133040, 32'sd1125312, 32'sd756457, 32'sd1113895, 32'sd1073546, 32'sd937936, 32'sd444372, 32'sd1038323,
32'sd791210, 32'sd954551, 32'sd502358, 32'sd997022, 32'sd1018741, 32'sd950310, 32'sd587189, 32'sd821419, 32'sd1150275, 32'sd1180292, 32'sd480688, 32'sd1160528, 32'sd829374, 32'sd1186080,
32'sd667806, 32'sd586205, 32'sd658856, 32'sd767503, 32'sd888459, 32'sd840204, 32'sd786232, 32'sd948674, 32'sd1151459, 32'sd1172207, 32'sd792207, 32'sd445473, 32'sd921736, 32'sd545531,
32'sd1201220, 32'sd785367, 32'sd603994, 32'sd779804, 32'sd580121, 32'sd634613, 32'sd731137, 32'sd437828, 32'sd1157278, 32'sd662025, 32'sd1012843, 32'sd934475, 32'sd688018, 32'sd1125817,
32'sd885753, 32'sd1114010, 32'sd1185787, 32'sd992658, 32'sd760169, 32'sd1060540, 32'sd824695, 32'sd994266, 32'sd459407, 32'sd1176442, 32'sd416779, 32'sd1039744, 32'sd440215, 32'sd1175494,
32'sd843290, 32'sd647330, 32'sd421987, 32'sd560844, 32'sd649745, 32'sd463697, 32'sd926359, 32'sd850595, 32'sd632993, 32'sd893762, 32'sd886916, 32'sd859701, 32'sd447271, 32'sd454883,
32'sd512038, 32'sd857700, 32'sd614567, 32'sd867810, 32'sd442490, 32'sd1133759, 32'sd865028, 32'sd878065, 32'sd645678, 32'sd471994, 32'sd643500, 32'sd1167289, 32'sd434260, 32'sd1196123,
32'sd824996, 32'sd864309, 32'sd446317, 32'sd924204, 32'sd462729, 32'sd917628, 32'sd581943, 32'sd646583, 32'sd817654, 32'sd605037, 32'sd1197369, 32'sd733001, 32'sd1206606, 32'sd769829,
32'sd1142787, 32'sd476878, 32'sd642196, 32'sd441439, 32'sd893835, 32'sd919170, 32'sd1182749, 32'sd658316, 32'sd831888, 32'sd1173207, 32'sd589073, 32'sd442189, 32'sd858256, 32'sd893172,
32'sd902220, 32'sd736562, 32'sd539250, 32'sd878741, 32'sd802703, 32'sd1138557, 32'sd1067284, 32'sd941298, 32'sd585386, 32'sd930694, 32'sd603006, 32'sd752907, 32'sd462010, 32'sd1012199,
32'sd409277, 32'sd1151614, 32'sd1003173, 32'sd617085, 32'sd1072931, 32'sd1136301, 32'sd650007, 32'sd635051, 32'sd519475, 32'sd1050256, 32'sd777544, 32'sd1046340, 32'sd1079199, 32'sd678491,
32'sd519985, 32'sd1184128, 32'sd497025, 32'sd907139, 32'sd911230, 32'sd1195053, 32'sd933862, 32'sd811625, 32'sd570653, 32'sd715707, 32'sd1051423, 32'sd1093358, 32'sd529273, 32'sd1033258,
32'sd1197689, 32'sd1101333, 32'sd630528, 32'sd643253, 32'sd742785, 32'sd628512, 32'sd767990, 32'sd486421, 32'sd528451, 32'sd580024, 32'sd704623, 32'sd852020, 32'sd595169, 32'sd1168095,
32'sd975689, 32'sd563882, 32'sd1086972, 32'sd969981, 32'sd602709, 32'sd981409, 32'sd881839, 32'sd553789, 32'sd614577, 32'sd890186, 32'sd763470, 32'sd977266, 32'sd889464, 32'sd719179,
32'sd888127, 32'sd781729, 32'sd978704, 32'sd492142, 32'sd828038, 32'sd1134556, 32'sd698388, 32'sd1160259, 32'sd832537, 32'sd481149, 32'sd888076, 32'sd624074, 32'sd1058211, 32'sd544433,
32'sd1018758, 32'sd754924, 32'sd1131745, 32'sd665976, 32'sd1125320, 32'sd856471, 32'sd558815, 32'sd807107, 32'sd524213, 32'sd662019, 32'sd1126563, 32'sd425977, 32'sd1089798, 32'sd1048113,
32'sd661819, 32'sd760560, 32'sd525396, 32'sd1135659, 32'sd707590, 32'sd1161324, 32'sd822270, 32'sd440482, 32'sd575111, 32'sd1051651, 32'sd1153614, 32'sd584709, 32'sd641435, 32'sd1195349,
32'sd981863, 32'sd767124, 32'sd645739, 32'sd863256, 32'sd461958, 32'sd425324, 32'sd1154104, 32'sd1185354, 32'sd973893, 32'sd618041, 32'sd465638, 32'sd1020471, 32'sd874619, 32'sd1007605,
32'sd773761, 32'sd985810, 32'sd542517, 32'sd1129069, 32'sd537665, 32'sd1014000, 32'sd906827, 32'sd417553, 32'sd1185013, 32'sd1015051, 32'sd753818, 32'sd791437, 32'sd839730, 32'sd707501,
32'sd701321, 32'sd539064, 32'sd740143, 32'sd731613, 32'sd456289, 32'sd580004, 32'sd1144715, 32'sd1134616, 32'sd922812, 32'sd757512, 32'sd787613, 32'sd1206568, 32'sd591826, 32'sd949698,
32'sd1021379, 32'sd573956, 32'sd1147538, 32'sd913502, 32'sd607045, 32'sd906236, 32'sd626493, 32'sd876818, 32'sd1005676, 32'sd561860, 32'sd1088591, 32'sd696363, 32'sd1134820, 32'sd1081097,
32'sd1031596, 32'sd737335, 32'sd716080, 32'sd514073, 32'sd919920, 32'sd511820, 32'sd966536, 32'sd434090, 32'sd885206, 32'sd524903, 32'sd746766, 32'sd1029423, 32'sd448965, 32'sd910766,
32'sd1209564, 32'sd548175, 32'sd512433, 32'sd601160, 32'sd979064, 32'sd862131, 32'sd894640, 32'sd679341, 32'sd1184742, 32'sd583661, 32'sd1144794, 32'sd1159396, 32'sd456134, 32'sd442448,
32'sd496779, 32'sd511394, 32'sd905245, 32'sd442909, 32'sd509815, 32'sd925744, 32'sd971750, 32'sd623930, 32'sd469584, 32'sd423442, 32'sd1031923, 32'sd706069, 32'sd1149375, 32'sd1142352,
32'sd1113863, 32'sd469024, 32'sd1042349, 32'sd949610, 32'sd926992, 32'sd1131646, 32'sd630105, 32'sd1030656, 32'sd1148513, 32'sd1198264, 32'sd753858, 32'sd970550, 32'sd522306, 32'sd923171,
32'sd722634, 32'sd1150568, 32'sd968604, 32'sd704460, 32'sd760408, 32'sd905035, 32'sd1050684, 32'sd1030003, 32'sd779695, 32'sd716217, 32'sd1051038, 32'sd701296, 32'sd568086, 32'sd1107531,
32'sd515558, 32'sd940989, 32'sd1044775, 32'sd476346, 32'sd827629, 32'sd707125, 32'sd648951, 32'sd507980, 32'sd1062141, 32'sd656283, 32'sd542175, 32'sd582825, 32'sd481438, 32'sd673285,
32'sd529147, 32'sd1184811, 32'sd518587, 32'sd1152889, 32'sd1171593, 32'sd915507, 32'sd805634, 32'sd961974, 32'sd441750, 32'sd1202753, 32'sd442913, 32'sd457209, 32'sd970190, 32'sd1123325,
32'sd998197, 32'sd689887, 32'sd1026109, 32'sd818114, 32'sd473552, 32'sd1091517, 32'sd677624, 32'sd908785, 32'sd656231, 32'sd484215, 32'sd1067162, 32'sd1103361, 32'sd1117191, 32'sd918249,
32'sd597633, 32'sd1204672, 32'sd507270, 32'sd802582, 32'sd632605, 32'sd1204741, 32'sd1089779, 32'sd501078, 32'sd1159749, 32'sd869597, 32'sd917767, 32'sd570509, 32'sd673933, 32'sd1093627,
32'sd824464, 32'sd910769, 32'sd1008480, 32'sd1137216, 32'sd1079182, 32'sd785165, 32'sd514121, 32'sd912770, 32'sd882937, 32'sd1150949, 32'sd820475, 32'sd817254, 32'sd826063, 32'sd731849,
32'sd431416, 32'sd1125762, 32'sd735246, 32'sd889245, 32'sd1076805, 32'sd700705, 32'sd862389, 32'sd1205014, 32'sd1148598, 32'sd823343, 32'sd787730, 32'sd796384, 32'sd938123, 32'sd1157515,
32'sd1117236, 32'sd1112244, 32'sd436063, 32'sd1100953, 32'sd500339, 32'sd772420, 32'sd788465, 32'sd502480, 32'sd638475, 32'sd801863, 32'sd712620, 32'sd823878, 32'sd412070, 32'sd832915,
32'sd884995, 32'sd484151, 32'sd1209171, 32'sd786094, 32'sd581725, 32'sd1123612, 32'sd669286, 32'sd457575, 32'sd452807, 32'sd690456, 32'sd867595, 32'sd779177, 32'sd449591, 32'sd567100,
32'sd693859, 32'sd553883, 32'sd449560, 32'sd871794, 32'sd858096, 32'sd906322, 32'sd905911, 32'sd837509, 32'sd407224, 32'sd1164596, 32'sd1077010, 32'sd1044093, 32'sd601928, 32'sd930649,
32'sd579186, 32'sd417511, 32'sd567172, 32'sd967280, 32'sd848637, 32'sd410765, 32'sd1185608, 32'sd1123084, 32'sd1206347, 32'sd481785, 32'sd1184278, 32'sd610130, 32'sd934312, 32'sd667576,
32'sd895688, 32'sd958833, 32'sd628635, 32'sd1073280, 32'sd588427, 32'sd1182789, 32'sd537754, 32'sd858062, 32'sd712777, 32'sd541874, 32'sd729028, 32'sd438740, 32'sd706903, 32'sd1202170,
32'sd550112, 32'sd648647, 32'sd1059441, 32'sd887132, 32'sd830742, 32'sd827350, 32'sd1135364, 32'sd409990, 32'sd908561, 32'sd764065, 32'sd557080, 32'sd572227, 32'sd1127882, 32'sd794179,
32'sd886085, 32'sd528585, 32'sd836381, 32'sd915817, 32'sd1007370, 32'sd1146584, 32'sd534217, 32'sd589368, 32'sd426203, 32'sd577467, 32'sd1179253, 32'sd1145060, 32'sd431378, 32'sd565657,
32'sd431311, 32'sd458870, 32'sd1173392, 32'sd1207021, 32'sd729186, 32'sd777657, 32'sd433912, 32'sd475597, 32'sd1042276, 32'sd1006995, 32'sd511964, 32'sd1183231, 32'sd578582, 32'sd1116567,
32'sd1047402, 32'sd884071, 32'sd823384, 32'sd629355, 32'sd556277, 32'sd697730, 32'sd885866, 32'sd1041795, 32'sd566817, 32'sd1103224, 32'sd1186676, 32'sd906140, 32'sd1034017, 32'sd511980,
32'sd1207195, 32'sd956441, 32'sd1140208, 32'sd755735, 32'sd1072653, 32'sd538023, 32'sd410521, 32'sd969956, 32'sd966310, 32'sd948169, 32'sd788643, 32'sd1081498, 32'sd679741, 32'sd969879,
32'sd1172733, 32'sd457153, 32'sd411370, 32'sd666162, 32'sd658865, 32'sd1189077, 32'sd1025334, 32'sd458332, 32'sd656316, 32'sd577183, 32'sd441694, 32'sd987560, 32'sd785393, 32'sd1049121,
32'sd1126734, 32'sd515760, 32'sd725650, 32'sd1054092, 32'sd1006996, 32'sd831443, 32'sd1188665, 32'sd920371, 32'sd956921, 32'sd819312, 32'sd685277, 32'sd555949, 32'sd424397, 32'sd720909,
32'sd475281, 32'sd515813, 32'sd722690, 32'sd884971, 32'sd489218, 32'sd845305, 32'sd926565, 32'sd636090, 32'sd783581, 32'sd449025, 32'sd798480, 32'sd1160076, 32'sd800989, 32'sd1012585,
32'sd902924, 32'sd857074, 32'sd1112054, 32'sd1154792, 32'sd524482, 32'sd1209063, 32'sd1015646, 32'sd506586, 32'sd1097396, 32'sd702851, 32'sd691124, 32'sd858269, 32'sd770511, 32'sd906468,
32'sd650827, 32'sd793717, 32'sd413935, 32'sd680534, 32'sd656149, 32'sd838903, 32'sd865352, 32'sd909508, 32'sd573231, 32'sd1140216, 32'sd496436, 32'sd482333, 32'sd1011775, 32'sd658022,
32'sd631747, 32'sd665040, 32'sd649094, 32'sd976966, 32'sd912469, 32'sd694431, 32'sd716506, 32'sd897719, 32'sd774116, 32'sd828013, 32'sd1092699, 32'sd1120710, 32'sd800913, 32'sd651414,
32'sd990968, 32'sd854677, 32'sd521439, 32'sd779174, 32'sd588832, 32'sd610323, 32'sd1048769, 32'sd451856, 32'sd1138910, 32'sd435181, 32'sd608131, 32'sd752414, 32'sd823132, 32'sd1202815,
32'sd842519, 32'sd969452, 32'sd826734, 32'sd771565, 32'sd709622, 32'sd782999, 32'sd456617, 32'sd928016, 32'sd1077922, 32'sd1095144, 32'sd903052, 32'sd838530, 32'sd736412, 32'sd1187568,
32'sd1200023, 32'sd1091272, 32'sd502340, 32'sd943997, 32'sd661098, 32'sd1017083, 32'sd1124232, 32'sd1109341, 32'sd859193, 32'sd1009167, 32'sd475185, 32'sd647000, 32'sd1171349, 32'sd561891,
32'sd693178, 32'sd408329, 32'sd560390, 32'sd902493, 32'sd494633, 32'sd782746, 32'sd660247, 32'sd964030, 32'sd844960, 32'sd1027109, 32'sd993320, 32'sd517931, 32'sd1050563, 32'sd653713,
32'sd895275, 32'sd1080938, 32'sd1117818, 32'sd404439, 32'sd689603, 32'sd1092816, 32'sd1175250, 32'sd552312, 32'sd938992, 32'sd848748, 32'sd945910, 32'sd715829, 32'sd715010, 32'sd482400,
32'sd969026, 32'sd984040, 32'sd690273, 32'sd1016928, 32'sd1130052, 32'sd921930, 32'sd866974, 32'sd918882, 32'sd957562, 32'sd1192716, 32'sd553805, 32'sd742663, 32'sd1179251, 32'sd855991,
32'sd758856, 32'sd612386, 32'sd1063818, 32'sd1070592, 32'sd550879, 32'sd859263, 32'sd902590, 32'sd1066916, 32'sd624121, 32'sd881296, 32'sd555528, 32'sd876331, 32'sd866960, 32'sd1001995,
32'sd881237, 32'sd457684, 32'sd861228, 32'sd502621, 32'sd1065592, 32'sd1181959, 32'sd1066741, 32'sd503214, 32'sd638995, 32'sd1130457, 32'sd575318, 32'sd418421, 32'sd1054061, 32'sd969643,
32'sd922342, 32'sd730669, 32'sd1155704, 32'sd1077068, 32'sd874721, 32'sd1016039, 32'sd776678, 32'sd1133643, 32'sd768061, 32'sd1039058, 32'sd814805, 32'sd989047, 32'sd852248, 32'sd1032931,
32'sd441535, 32'sd784679, 32'sd652299, 32'sd1033780, 32'sd556238, 32'sd776922, 32'sd1030832, 32'sd837814, 32'sd1087113, 32'sd1066758, 32'sd1156553, 32'sd730122, 32'sd864230, 32'sd616454,
32'sd597253, 32'sd573504, 32'sd1023864, 32'sd800845, 32'sd739365, 32'sd1080532, 32'sd461209, 32'sd829761, 32'sd568873, 32'sd1103587, 32'sd420897, 32'sd1052879, 32'sd484973, 32'sd1096459,
32'sd790402, 32'sd458648, 32'sd430251, 32'sd782501, 32'sd550390, 32'sd1164443, 32'sd1104533, 32'sd697075, 32'sd619724, 32'sd800017, 32'sd891971, 32'sd1200244, 32'sd429376, 32'sd649417,
32'sd586265, 32'sd557355, 32'sd864464, 32'sd803742, 32'sd644940, 32'sd1111842, 32'sd636017, 32'sd603736, 32'sd485064, 32'sd781539, 32'sd869459, 32'sd635386, 32'sd712835, 32'sd1020625,
32'sd756331, 32'sd1178811, 32'sd1081645, 32'sd829629, 32'sd818344, 32'sd1074290, 32'sd913332, 32'sd679801, 32'sd990214, 32'sd474536, 32'sd904732, 32'sd1137012, 32'sd850605, 32'sd1162865,
32'sd1021016, 32'sd1028507, 32'sd929594, 32'sd432609, 32'sd991275, 32'sd834908, 32'sd924542, 32'sd544457, 32'sd1204731, 32'sd660874, 32'sd826717, 32'sd677376, 32'sd1118643, 32'sd568394,
32'sd919180, 32'sd930460, 32'sd492208, 32'sd914098, 32'sd698122, 32'sd1008080, 32'sd529523, 32'sd545119, 32'sd591697, 32'sd624754, 32'sd1022415, 32'sd952856, 32'sd940240, 32'sd959581,
32'sd1134616, 32'sd996105, 32'sd958462, 32'sd649730, 32'sd812631, 32'sd884835, 32'sd981588, 32'sd699407, 32'sd616515, 32'sd1177407, 32'sd681985, 32'sd1013941, 32'sd1159981, 32'sd622265,
32'sd422000, 32'sd453233, 32'sd556906, 32'sd972446, 32'sd606390, 32'sd518734, 32'sd937598, 32'sd862685, 32'sd1082917, 32'sd675178, 32'sd1142166, 32'sd850721, 32'sd799317, 32'sd674229,
32'sd804130, 32'sd748256, 32'sd669396, 32'sd490562, 32'sd612378, 32'sd851158, 32'sd887576, 32'sd511071, 32'sd992604, 32'sd1103679, 32'sd1154548, 32'sd1188949, 32'sd597482, 32'sd1088962,
32'sd1149105, 32'sd968061, 32'sd654164, 32'sd597818, 32'sd414831, 32'sd987736, 32'sd1205658, 32'sd966630, 32'sd944102, 32'sd507521, 32'sd786878, 32'sd1119568, 32'sd895768, 32'sd479429,
32'sd795622, 32'sd588067, 32'sd648421, 32'sd1115214, 32'sd787982, 32'sd767809, 32'sd956455, 32'sd1057826, 32'sd813277, 32'sd975903, 32'sd502120, 32'sd1161535, 32'sd745901, 32'sd661752,
32'sd866727, 32'sd1025226, 32'sd486972, 32'sd855280, 32'sd671675, 32'sd1142613, 32'sd1076529, 32'sd743508, 32'sd646000, 32'sd823144, 32'sd444345, 32'sd578408, 32'sd547724, 32'sd728575,
32'sd847857, 32'sd984820, 32'sd963679, 32'sd619752, 32'sd471981, 32'sd606261, 32'sd419364, 32'sd597526, 32'sd473231, 32'sd979720, 32'sd1168335, 32'sd804426, 32'sd768101, 32'sd769460,
32'sd880042, 32'sd678931, 32'sd499364, 32'sd459113, 32'sd716514, 32'sd1111206, 32'sd590733, 32'sd577006, 32'sd649386, 32'sd1126311, 32'sd525053, 32'sd1053497, 32'sd681283, 32'sd872598,
32'sd592364, 32'sd884862, 32'sd672670, 32'sd1168145, 32'sd1185951, 32'sd869430, 32'sd492474, 32'sd506925, 32'sd462150, 32'sd673697, 32'sd898838, 32'sd887555, 32'sd753302, 32'sd914915,
32'sd467350, 32'sd822661, 32'sd544076, 32'sd780046, 32'sd621958, 32'sd411557, 32'sd557192, 32'sd721369, 32'sd542252, 32'sd1007651, 32'sd531883, 32'sd916580, 32'sd485997, 32'sd539460,
32'sd897851, 32'sd550902, 32'sd1105137, 32'sd941438, 32'sd1192424, 32'sd1184866, 32'sd1135461, 32'sd783669, 32'sd662223, 32'sd549346, 32'sd456275, 32'sd583324, 32'sd552969, 32'sd871954,
32'sd598798, 32'sd982064, 32'sd886497, 32'sd1188576, 32'sd689816, 32'sd532483, 32'sd426923, 32'sd547954, 32'sd679514, 32'sd558638, 32'sd904554, 32'sd995126, 32'sd1146821, 32'sd751348,
32'sd536508, 32'sd791328, 32'sd754220, 32'sd808110, 32'sd694187, 32'sd989506, 32'sd781775, 32'sd812144, 32'sd616109, 32'sd550921, 32'sd777524, 32'sd677321, 32'sd582884, 32'sd973372,
32'sd994363, 32'sd951836, 32'sd423478, 32'sd432651, 32'sd603508, 32'sd548901, 32'sd1173348, 32'sd843480, 32'sd610288, 32'sd949663, 32'sd1138870, 32'sd459875, 32'sd592637, 32'sd1073713,
32'sd767878, 32'sd989946, 32'sd579276, 32'sd1139413, 32'sd974951, 32'sd1060257, 32'sd998565, 32'sd785504, 32'sd537137, 32'sd926838, 32'sd439071, 32'sd792670, 32'sd1141275, 32'sd1084999,
32'sd405310, 32'sd861816, 32'sd577885, 32'sd408363, 32'sd851427, 32'sd744582, 32'sd1035361, 32'sd747878, 32'sd424038, 32'sd1114657, 32'sd912449, 32'sd744129, 32'sd979391, 32'sd954119,
32'sd565234, 32'sd549110, 32'sd1180449, 32'sd647318, 32'sd560258, 32'sd1130845, 32'sd930181, 32'sd926460, 32'sd465353, 32'sd1101796, 32'sd772163, 32'sd1052668, 32'sd1093476, 32'sd631426,
32'sd667266, 32'sd1165196, 32'sd496736, 32'sd414795, 32'sd916670, 32'sd681277, 32'sd710306, 32'sd462973, 32'sd580179, 32'sd470804, 32'sd1204791, 32'sd1162603, 32'sd983890, 32'sd1067321,
32'sd590364, 32'sd1189675, 32'sd510390, 32'sd408217, 32'sd1111138, 32'sd1155917, 32'sd1045602, 32'sd727947, 32'sd738900, 32'sd801468, 32'sd564851, 32'sd1178198, 32'sd596009, 32'sd1112242,
32'sd1007839, 32'sd684691, 32'sd985209, 32'sd795349, 32'sd1030695, 32'sd812107, 32'sd917744, 32'sd1110928, 32'sd1034069, 32'sd819404, 32'sd665923, 32'sd794783, 32'sd1140128, 32'sd859595,
32'sd572418, 32'sd916863, 32'sd1149387, 32'sd1057891, 32'sd681132, 32'sd447415, 32'sd913862, 32'sd779447, 32'sd1167559, 32'sd1205834, 32'sd676508, 32'sd1073907, 32'sd1205577, 32'sd585115,
32'sd755002, 32'sd873898, 32'sd1129091, 32'sd613537, 32'sd415260, 32'sd625879, 32'sd494931, 32'sd415756, 32'sd921433, 32'sd1129681, 32'sd591238, 32'sd696496, 32'sd638777, 32'sd908947,
32'sd854673, 32'sd1056097, 32'sd415833, 32'sd475231, 32'sd1201892, 32'sd919668, 32'sd457316, 32'sd600937, 32'sd746647, 32'sd414658, 32'sd967691, 32'sd629822, 32'sd995976, 32'sd664130,
32'sd418399, 32'sd928906, 32'sd865422, 32'sd1070386, 32'sd1160387, 32'sd920717, 32'sd409643, 32'sd491789, 32'sd562565, 32'sd505672, 32'sd758892, 32'sd704399, 32'sd1170356, 32'sd534427,
32'sd461728, 32'sd864792, 32'sd812646, 32'sd1055353, 32'sd906835, 32'sd874916, 32'sd403847, 32'sd874499, 32'sd428871, 32'sd627229, 32'sd897465, 32'sd889845, 32'sd629604, 32'sd810835,
32'sd1132812, 32'sd822077, 32'sd491375, 32'sd928660, 32'sd531074, 32'sd841329, 32'sd429511, 32'sd1175129, 32'sd687042, 32'sd553639, 32'sd834571, 32'sd655221, 32'sd759668, 32'sd522902,
32'sd699224, 32'sd543987, 32'sd1095192, 32'sd732550, 32'sd873723, 32'sd1038137, 32'sd503322, 32'sd980674, 32'sd1135815, 32'sd1008257, 32'sd472886, 32'sd836837, 32'sd458103, 32'sd1203218,
32'sd1140157, 32'sd437763, 32'sd572562, 32'sd845900, 32'sd473780, 32'sd442590, 32'sd925896, 32'sd803749, 32'sd451352, 32'sd601253, 32'sd985143, 32'sd715723, 32'sd531214, 32'sd807403,
32'sd517973, 32'sd671165, 32'sd779209, 32'sd475220, 32'sd1076183, 32'sd1083299, 32'sd692037, 32'sd570181, 32'sd601731, 32'sd433366, 32'sd659993, 32'sd926513, 32'sd1197852, 32'sd784797,
32'sd677360, 32'sd426256, 32'sd451507, 32'sd1104887, 32'sd605021, 32'sd1015568, 32'sd519710, 32'sd661392, 32'sd572163, 32'sd826351, 32'sd698894, 32'sd681809, 32'sd1091524, 32'sd719321,
32'sd544996, 32'sd746484, 32'sd1193921, 32'sd613305, 32'sd1071692, 32'sd1076178, 32'sd598474, 32'sd968270, 32'sd894343, 32'sd1014657, 32'sd747089, 32'sd939013, 32'sd993351, 32'sd857355,
32'sd990527, 32'sd1037225, 32'sd616747, 32'sd1183666, 32'sd895035, 32'sd963533, 32'sd477006, 32'sd754554, 32'sd665390, 32'sd904579, 32'sd1180475, 32'sd481610, 32'sd937146, 32'sd858145,
32'sd768736, 32'sd626399, 32'sd966505, 32'sd468543, 32'sd523987, 32'sd538263, 32'sd1024256, 32'sd1164534, 32'sd483214, 32'sd429808, 32'sd707401, 32'sd1082487, 32'sd906608, 32'sd902064,
32'sd712453, 32'sd1191121, 32'sd691844, 32'sd1091449, 32'sd739847, 32'sd908045, 32'sd756027, 32'sd460499, 32'sd1170637, 32'sd588445, 32'sd978686, 32'sd614319, 32'sd1170888, 32'sd1111386,
32'sd966824, 32'sd1038796, 32'sd561265, 32'sd784147, 32'sd664663, 32'sd1026587, 32'sd457971, 32'sd1060332, 32'sd912592, 32'sd443384, 32'sd790860, 32'sd510059, 32'sd818094, 32'sd1115656,
32'sd503224, 32'sd631199, 32'sd978178, 32'sd1067761, 32'sd664525, 32'sd504543, 32'sd904921, 32'sd881917, 32'sd609339, 32'sd1067995, 32'sd662532, 32'sd761164, 32'sd1084677, 32'sd565158,
32'sd490445, 32'sd1029506, 32'sd947940, 32'sd1154435, 32'sd1149757, 32'sd792058, 32'sd590927, 32'sd1134092, 32'sd924215, 32'sd557991, 32'sd949852, 32'sd648192, 32'sd677594, 32'sd915341,
32'sd634949, 32'sd1156930, 32'sd549050, 32'sd1045110, 32'sd555357, 32'sd704750, 32'sd584220, 32'sd851710, 32'sd684934, 32'sd1029034, 32'sd472015, 32'sd772195, 32'sd898050, 32'sd541678,
32'sd1059477, 32'sd979650, 32'sd1131206, 32'sd416303, 32'sd1132006, 32'sd722161, 32'sd1096250, 32'sd521591, 32'sd923808, 32'sd713442, 32'sd939508, 32'sd1137352, 32'sd991062, 32'sd895508,
32'sd559887, 32'sd801345, 32'sd542476, 32'sd1102304, 32'sd794129, 32'sd1009549, 32'sd1057993, 32'sd711065, 32'sd859907, 32'sd1120908, 32'sd538037, 32'sd948023, 32'sd495872, 32'sd851462,
32'sd1100072, 32'sd696060, 32'sd610281, 32'sd924181, 32'sd535806, 32'sd709209, 32'sd446689, 32'sd1010568, 32'sd780102, 32'sd570711, 32'sd760201, 32'sd752256, 32'sd951401, 32'sd794295,
32'sd588696, 32'sd979120, 32'sd1171071, 32'sd880041, 32'sd764965, 32'sd681010, 32'sd978224, 32'sd953239, 32'sd919114, 32'sd1056719, 32'sd916394, 32'sd755311, 32'sd882475, 32'sd504404,
32'sd1002900, 32'sd792067, 32'sd1199141, 32'sd688960, 32'sd1027870, 32'sd897510, 32'sd724178, 32'sd989992, 32'sd752841, 32'sd614826, 32'sd727010, 32'sd676650, 32'sd1061707, 32'sd1150907,
32'sd521001, 32'sd1053883, 32'sd777403, 32'sd1099553, 32'sd1076126, 32'sd567571, 32'sd896221, 32'sd653298, 32'sd987231, 32'sd1192858, 32'sd1139783, 32'sd839851, 32'sd1202341, 32'sd1155662,
32'sd628303, 32'sd760194, 32'sd723385, 32'sd475610, 32'sd658960, 32'sd1147326, 32'sd947186, 32'sd1084533, 32'sd554842, 32'sd992498, 32'sd610199, 32'sd1125443, 32'sd547563, 32'sd683313,
32'sd546578, 32'sd465433, 32'sd937868, 32'sd1174234, 32'sd758272, 32'sd529035, 32'sd972768, 32'sd419313, 32'sd657308, 32'sd784162, 32'sd1095557, 32'sd960255, 32'sd1141108, 32'sd765347,
32'sd703828, 32'sd869167, 32'sd1063975, 32'sd915251, 32'sd550402, 32'sd660629, 32'sd978374, 32'sd786003, 32'sd1079954, 32'sd976436, 32'sd478162, 32'sd606591, 32'sd1161612, 32'sd407730,
32'sd1029236, 32'sd569756, 32'sd787550, 32'sd460881, 32'sd1032852, 32'sd540904, 32'sd853650, 32'sd1026042, 32'sd428555, 32'sd659478, 32'sd789546, 32'sd1096592, 32'sd958237, 32'sd438398,
32'sd573442, 32'sd970191, 32'sd460498, 32'sd788222, 32'sd901368, 32'sd898421, 32'sd897691, 32'sd542827, 32'sd557759, 32'sd820454, 32'sd483595, 32'sd1171117, 32'sd808667, 32'sd1069953,
32'sd605236, 32'sd951065, 32'sd439162, 32'sd1105185, 32'sd655356, 32'sd596405, 32'sd982617, 32'sd796761, 32'sd845515, 32'sd1113438, 32'sd1130390, 32'sd566690, 32'sd804480, 32'sd799751,
32'sd1064639, 32'sd722337, 32'sd806410, 32'sd979815, 32'sd459649, 32'sd858289, 32'sd773765, 32'sd942362, 32'sd922252, 32'sd1094400, 32'sd1103389, 32'sd460213, 32'sd874500, 32'sd532159,
32'sd650482, 32'sd837838, 32'sd1086826, 32'sd970229, 32'sd863709, 32'sd488732, 32'sd1085573, 32'sd938200, 32'sd951717, 32'sd444364, 32'sd1167196, 32'sd1010926, 32'sd964537, 32'sd882004,
32'sd540340, 32'sd464322, 32'sd1209099, 32'sd521054, 32'sd1112503, 32'sd818918, 32'sd494857, 32'sd686933, 32'sd813192, 32'sd604775, 32'sd1153762, 32'sd915988, 32'sd928305, 32'sd751535,
32'sd957719, 32'sd524147, 32'sd1082076, 32'sd1084266, 32'sd928612, 32'sd549684, 32'sd896910, 32'sd1134177, 32'sd494338, 32'sd809677, 32'sd1129335, 32'sd790564, 32'sd689581, 32'sd1199995,
32'sd754046, 32'sd916798, 32'sd1132836, 32'sd773291, 32'sd1154113, 32'sd522438, 32'sd436003, 32'sd1022020, 32'sd426227, 32'sd1095644, 32'sd925762, 32'sd804207, 32'sd791813, 32'sd992913,
32'sd551297, 32'sd671722, 32'sd577268, 32'sd1152555, 32'sd1018551, 32'sd494448, 32'sd405984, 32'sd1147602, 32'sd582486, 32'sd673026, 32'sd867711, 32'sd820521, 32'sd737976, 32'sd629716,
32'sd657075, 32'sd773292, 32'sd527911, 32'sd861422, 32'sd740524, 32'sd604216, 32'sd527181, 32'sd1007225, 32'sd921931, 32'sd885523, 32'sd561052, 32'sd1174127, 32'sd1048666, 32'sd410269,
32'sd803740, 32'sd862623, 32'sd848136, 32'sd977499, 32'sd616628, 32'sd910940, 32'sd1114043, 32'sd1073888, 32'sd505633, 32'sd1134212, 32'sd739950, 32'sd683702, 32'sd1090799, 32'sd817761,
32'sd789472, 32'sd1094150, 32'sd1089659, 32'sd1060936, 32'sd799045, 32'sd610858, 32'sd1181531, 32'sd976065, 32'sd600102, 32'sd1187046, 32'sd924984, 32'sd532223, 32'sd466012, 32'sd1207541,
32'sd949083, 32'sd558429, 32'sd777170, 32'sd474078, 32'sd673118, 32'sd1057056, 32'sd1142599, 32'sd983725, 32'sd1179640, 32'sd1138605, 32'sd920785, 32'sd521999, 32'sd556323, 32'sd407082,
32'sd816071, 32'sd988795, 32'sd1156943, 32'sd754067, 32'sd704979, 32'sd1012185, 32'sd592733, 32'sd1041390, 32'sd772713, 32'sd840029, 32'sd1128134, 32'sd1200531, 32'sd936350, 32'sd1093646,
32'sd1076230, 32'sd750648, 32'sd826718, 32'sd1052002, 32'sd660811, 32'sd727727, 32'sd741523, 32'sd610307, 32'sd636435, 32'sd1006548, 32'sd785617, 32'sd688424, 32'sd1027602, 32'sd809433,
32'sd767075, 32'sd690668, 32'sd712921, 32'sd992576, 32'sd506780, 32'sd947162, 32'sd660003, 32'sd669874, 32'sd821625, 32'sd1046844, 32'sd1104885, 32'sd1141237, 32'sd561465, 32'sd562025,
32'sd440390, 32'sd948783, 32'sd428252, 32'sd914524, 32'sd1180432, 32'sd1198992, 32'sd735458, 32'sd676095, 32'sd679392, 32'sd1039053, 32'sd1098083, 32'sd682372, 32'sd881436, 32'sd650752,
32'sd735644, 32'sd540063, 32'sd831159, 32'sd1077280, 32'sd1075910, 32'sd980455, 32'sd491335, 32'sd1034348, 32'sd1163191, 32'sd1163479, 32'sd482153, 32'sd959990, 32'sd1079581, 32'sd839143,
32'sd905487, 32'sd945399, 32'sd778259, 32'sd479695, 32'sd405996, 32'sd752068, 32'sd962535, 32'sd564143, 32'sd1036672, 32'sd590748, 32'sd607025, 32'sd978147, 32'sd871937, 32'sd737965,
32'sd1142621, 32'sd905630, 32'sd1067995, 32'sd1040514, 32'sd658531, 32'sd565192, 32'sd701026, 32'sd837791, 32'sd896340, 32'sd974415, 32'sd601610, 32'sd1199024, 32'sd957189, 32'sd652963,
32'sd987487, 32'sd657148, 32'sd1051979, 32'sd1000553, 32'sd1049480, 32'sd733172, 32'sd1008854, 32'sd1053837, 32'sd915836, 32'sd1057580, 32'sd998133, 32'sd1198511, 32'sd601345, 32'sd1096675,
32'sd866765, 32'sd1118663, 32'sd1163699, 32'sd1179424, 32'sd1061543, 32'sd460717, 32'sd891997, 32'sd613107, 32'sd1057654, 32'sd900669, 32'sd994443, 32'sd1134460, 32'sd589423, 32'sd623859,
32'sd821684, 32'sd780846, 32'sd697481, 32'sd779178, 32'sd796446, 32'sd1168634, 32'sd462319, 32'sd887935, 32'sd901375, 32'sd980285, 32'sd561720, 32'sd930030, 32'sd570894, 32'sd791935,
32'sd761562, 32'sd730331, 32'sd793096, 32'sd823901, 32'sd1056847, 32'sd711949, 32'sd882913, 32'sd798451, 32'sd777536, 32'sd554943, 32'sd670679, 32'sd512983, 32'sd701847, 32'sd531724,
32'sd635725, 32'sd804911, 32'sd1072561, 32'sd998674, 32'sd812207, 32'sd1005362, 32'sd417622, 32'sd896375, 32'sd607129, 32'sd609922, 32'sd891563, 32'sd731160, 32'sd615374, 32'sd1036654,
32'sd503639, 32'sd500793, 32'sd680412, 32'sd789530, 32'sd498353, 32'sd1057535, 32'sd914070, 32'sd708212, 32'sd1059598, 32'sd878045, 32'sd501591, 32'sd643358, 32'sd610670, 32'sd521736,
32'sd544049, 32'sd1089696, 32'sd768138, 32'sd658834, 32'sd483945, 32'sd770342, 32'sd675988, 32'sd767542, 32'sd1075824, 32'sd1024308, 32'sd1013130, 32'sd988698, 32'sd1172433, 32'sd599687,
32'sd643077, 32'sd813655, 32'sd1034378, 32'sd823160, 32'sd1014353, 32'sd658349, 32'sd637057, 32'sd548884, 32'sd484961, 32'sd854544, 32'sd703476, 32'sd886282, 32'sd926282, 32'sd426261,
32'sd1175542, 32'sd606423, 32'sd1007229, 32'sd782517, 32'sd940519, 32'sd430408, 32'sd754162, 32'sd455359, 32'sd900558, 32'sd661279, 32'sd590217, 32'sd1070101, 32'sd587578, 32'sd624719,
32'sd638544, 32'sd1038799, 32'sd837896, 32'sd1023682, 32'sd686353, 32'sd766110, 32'sd625271, 32'sd430426, 32'sd495014, 32'sd630023, 32'sd866745, 32'sd743457, 32'sd1028095, 32'sd754049,
32'sd627372, 32'sd972341, 32'sd1080049, 32'sd489439, 32'sd605279, 32'sd1007917, 32'sd632264, 32'sd1110132, 32'sd775165, 32'sd728423, 32'sd660380, 32'sd497275, 32'sd816244, 32'sd710821,
32'sd806618, 32'sd488493, 32'sd1126159, 32'sd404775, 32'sd735919, 32'sd673330, 32'sd503312, 32'sd952364, 32'sd1156298, 32'sd1135071, 32'sd798333, 32'sd588534, 32'sd689300, 32'sd419711,
32'sd486409, 32'sd735848, 32'sd668786, 32'sd428452, 32'sd838935, 32'sd834137, 32'sd862244, 32'sd1128641, 32'sd952102, 32'sd1064748, 32'sd640286, 32'sd1018943, 32'sd471706, 32'sd1116446,
32'sd899807, 32'sd505397, 32'sd667967, 32'sd975021, 32'sd1057416, 32'sd1199539, 32'sd1063002, 32'sd867087, 32'sd1158305, 32'sd1177797, 32'sd403465, 32'sd1033841, 32'sd1144604, 32'sd1010137,
32'sd858076, 32'sd441784, 32'sd957192, 32'sd551062, 32'sd482309, 32'sd1205305, 32'sd1084622, 32'sd1174255, 32'sd536277, 32'sd1122661, 32'sd488805, 32'sd880053, 32'sd758109, 32'sd598240,
32'sd1091773, 32'sd1179474, 32'sd656557, 32'sd680522, 32'sd525552, 32'sd765019, 32'sd496832, 32'sd1199983, 32'sd756024, 32'sd639113, 32'sd694738, 32'sd1039422, 32'sd429221, 32'sd835557,
32'sd993934, 32'sd1120822, 32'sd858207, 32'sd885563, 32'sd865405, 32'sd847555, 32'sd787568, 32'sd815687, 32'sd468879, 32'sd994450, 32'sd981605, 32'sd1135584, 32'sd1139528, 32'sd1119273,
32'sd841620, 32'sd1108910, 32'sd1170450, 32'sd824813, 32'sd435503, 32'sd1098645, 32'sd903897, 32'sd667524, 32'sd1060170, 32'sd883419, 32'sd984677, 32'sd997730, 32'sd858304, 32'sd548181,
32'sd952979, 32'sd669262, 32'sd522275, 32'sd482579, 32'sd806019, 32'sd858550, 32'sd547626, 32'sd779216, 32'sd1057459, 32'sd788758, 32'sd1204041, 32'sd575883, 32'sd958365, 32'sd973090,
32'sd688279, 32'sd907971, 32'sd1129103, 32'sd708477, 32'sd433496, 32'sd1111858, 32'sd600136, 32'sd873290, 32'sd788832, 32'sd521685, 32'sd1150021, 32'sd909067, 32'sd752689, 32'sd599880,
32'sd708674, 32'sd1063333, 32'sd674359, 32'sd582061, 32'sd614142, 32'sd657857, 32'sd661231, 32'sd1084427, 32'sd791239, 32'sd998128, 32'sd524483, 32'sd1116197, 32'sd888852, 32'sd732878,
32'sd436221, 32'sd733359, 32'sd1186537, 32'sd1095973, 32'sd708995, 32'sd611016, 32'sd1041895, 32'sd590627, 32'sd738585, 32'sd586676, 32'sd558734, 32'sd529876, 32'sd485744, 32'sd904385,
32'sd596354, 32'sd878420, 32'sd1178088, 32'sd752410, 32'sd603111, 32'sd737819, 32'sd744054, 32'sd652844, 32'sd494094, 32'sd922253, 32'sd1110195, 32'sd990846, 32'sd1063850, 32'sd443427,
32'sd1207488, 32'sd605460, 32'sd633863, 32'sd459249, 32'sd1188026, 32'sd487415, 32'sd712204, 32'sd764288, 32'sd769177, 32'sd562123, 32'sd874055, 32'sd537318, 32'sd754658, 32'sd1115390,
32'sd1035052, 32'sd884423, 32'sd1165594, 32'sd1020914, 32'sd558573, 32'sd459469, 32'sd1150345, 32'sd1049636, 32'sd1149008, 32'sd1016102, 32'sd655371, 32'sd949401, 32'sd512275, 32'sd803315,
32'sd778050, 32'sd896654, 32'sd956458, 32'sd867305, 32'sd790764, 32'sd1163400, 32'sd892436, 32'sd653764, 32'sd867879, 32'sd1153659, 32'sd893947, 32'sd600204, 32'sd587570, 32'sd776814,
32'sd1059654, 32'sd494924, 32'sd703287, 32'sd802571, 32'sd1026216, 32'sd693145, 32'sd975668, 32'sd1054418, 32'sd986416, 32'sd805688, 32'sd695406, 32'sd540465, 32'sd1209383, 32'sd851429,
32'sd674536, 32'sd930737, 32'sd856060, 32'sd767749, 32'sd779421, 32'sd1170424, 32'sd622546, 32'sd501329, 32'sd494094, 32'sd1209157, 32'sd1000145, 32'sd772046, 32'sd1135929, 32'sd649752,
32'sd452274, 32'sd1138099, 32'sd598831, 32'sd444407, 32'sd1114392, 32'sd731218, 32'sd1058156, 32'sd857879, 32'sd853924, 32'sd906756, 32'sd518510, 32'sd982717, 32'sd640478, 32'sd1023640,
32'sd661972, 32'sd1157279, 32'sd583303, 32'sd468702, 32'sd610673, 32'sd1196587, 32'sd1057686, 32'sd1094984, 32'sd787015, 32'sd1006328, 32'sd679696, 32'sd901882, 32'sd588217, 32'sd645921,
32'sd1166007, 32'sd1077532, 32'sd1057777, 32'sd525009, 32'sd990187, 32'sd968927, 32'sd455805, 32'sd507927, 32'sd768703, 32'sd851530, 32'sd655087, 32'sd567066, 32'sd1166113, 32'sd1207828,
32'sd875649, 32'sd446896, 32'sd645336, 32'sd893777, 32'sd614425, 32'sd1082660, 32'sd810519, 32'sd441109, 32'sd1029470, 32'sd1020955, 32'sd906969, 32'sd1202585, 32'sd1062797, 32'sd576105,
32'sd487130, 32'sd607150, 32'sd621148, 32'sd719525, 32'sd638045, 32'sd982739, 32'sd1174588, 32'sd682800, 32'sd414787, 32'sd949636, 32'sd1149416, 32'sd446952, 32'sd646046, 32'sd1145206,
32'sd607004, 32'sd1201107, 32'sd508250, 32'sd1134901, 32'sd1066475, 32'sd533680, 32'sd943742, 32'sd758318, 32'sd586020, 32'sd453465, 32'sd1028376, 32'sd929405, 32'sd1088932, 32'sd1190911,
32'sd687743, 32'sd1026435, 32'sd910303, 32'sd827424, 32'sd767138, 32'sd734132, 32'sd1113950, 32'sd543085, 32'sd821729, 32'sd1104185, 32'sd1098700, 32'sd743397, 32'sd991423, 32'sd1034616,
32'sd911641, 32'sd906327, 32'sd1176355, 32'sd992877, 32'sd1099842, 32'sd860686, 32'sd946598, 32'sd704221, 32'sd812884, 32'sd993622, 32'sd1143409, 32'sd719785, 32'sd1031319, 32'sd1044036,
32'sd911204, 32'sd432798, 32'sd896102, 32'sd700940, 32'sd665209, 32'sd1168733, 32'sd1108983, 32'sd582077, 32'sd919841, 32'sd886942, 32'sd1068202, 32'sd484380, 32'sd1012942, 32'sd1082450,
32'sd541056, 32'sd775334, 32'sd1174792, 32'sd809307, 32'sd420026, 32'sd909484, 32'sd1007479, 32'sd862795, 32'sd1094504, 32'sd831151, 32'sd836938, 32'sd1148383, 32'sd500139, 32'sd1022372,
32'sd568526, 32'sd880669, 32'sd1151697, 32'sd850499, 32'sd1104986, 32'sd1085597, 32'sd1020778, 32'sd476425, 32'sd747528, 32'sd1058613, 32'sd443293, 32'sd872344, 32'sd663728, 32'sd1199208,
32'sd974299, 32'sd531503, 32'sd1071597, 32'sd1168266, 32'sd542554, 32'sd684332, 32'sd783532, 32'sd766359, 32'sd1207862, 32'sd1085692, 32'sd1141654, 32'sd945011, 32'sd723743, 32'sd725404,
32'sd693656, 32'sd845174, 32'sd451421, 32'sd411809, 32'sd734561, 32'sd420969, 32'sd579477, 32'sd819823, 32'sd668243, 32'sd491625, 32'sd653547, 32'sd475273, 32'sd473021, 32'sd870383,
32'sd590344, 32'sd456123, 32'sd727599, 32'sd1002087, 32'sd1179924, 32'sd643638, 32'sd834970, 32'sd836473, 32'sd1091584, 32'sd1016605, 32'sd1198355, 32'sd446130, 32'sd1026511, 32'sd1161798,
32'sd579002, 32'sd934737, 32'sd578939, 32'sd488131, 32'sd730383, 32'sd773132, 32'sd411390, 32'sd800517, 32'sd507492, 32'sd1073370, 32'sd1034458, 32'sd472301, 32'sd651096, 32'sd563953,
32'sd1021574, 32'sd719027, 32'sd1192166, 32'sd1205121, 32'sd959286, 32'sd1122842, 32'sd1080931, 32'sd1158916, 32'sd580083, 32'sd472727, 32'sd1034733, 32'sd473894, 32'sd1066793, 32'sd600882,
32'sd404867, 32'sd683714, 32'sd505938, 32'sd992260, 32'sd721514, 32'sd769474, 32'sd925452, 32'sd641184, 32'sd634937, 32'sd905654, 32'sd713660, 32'sd869837, 32'sd1126760, 32'sd1063542,
32'sd658586, 32'sd1182392, 32'sd594491, 32'sd1018940, 32'sd577895, 32'sd559652, 32'sd450775, 32'sd541057, 32'sd471539, 32'sd809780, 32'sd733383, 32'sd740941, 32'sd1163348, 32'sd483883,
32'sd567309, 32'sd634510, 32'sd1066883, 32'sd538807, 32'sd609775, 32'sd723790, 32'sd1128929, 32'sd928462, 32'sd1070103, 32'sd1143451, 32'sd938790, 32'sd1122011, 32'sd1129423, 32'sd1174349,
32'sd902404, 32'sd529754, 32'sd630472, 32'sd1130315, 32'sd1082845, 32'sd935454, 32'sd1068008, 32'sd851322, 32'sd434221, 32'sd657111, 32'sd709551, 32'sd572031, 32'sd919555, 32'sd775756,
32'sd891853, 32'sd1009933, 32'sd416448, 32'sd403556, 32'sd875736, 32'sd829818, 32'sd868098, 32'sd825963, 32'sd711511, 32'sd681706, 32'sd1177263, 32'sd456629, 32'sd676973, 32'sd888214,
32'sd624280, 32'sd915439, 32'sd707961, 32'sd687265, 32'sd405432, 32'sd929759, 32'sd1082301, 32'sd477213, 32'sd473264, 32'sd636810, 32'sd879447, 32'sd756738, 32'sd1195245, 32'sd642933,
32'sd466632, 32'sd738805, 32'sd560372, 32'sd426323, 32'sd566817, 32'sd626467, 32'sd476192, 32'sd609174, 32'sd549699, 32'sd841506, 32'sd720412, 32'sd871814, 32'sd924618, 32'sd753694,
32'sd950297, 32'sd474936, 32'sd522464, 32'sd947031, 32'sd636460, 32'sd1103538, 32'sd967444, 32'sd882041, 32'sd769953, 32'sd974374, 32'sd416381, 32'sd478812, 32'sd538684, 32'sd646857,
32'sd934795, 32'sd684214, 32'sd593731, 32'sd623871, 32'sd465749, 32'sd532826, 32'sd495258, 32'sd555244, 32'sd958355, 32'sd736487, 32'sd475309, 32'sd762063, 32'sd631014, 32'sd708862,
32'sd740621, 32'sd699065, 32'sd1197139, 32'sd746667, 32'sd1082452, 32'sd420914, 32'sd1189344, 32'sd979872, 32'sd592131, 32'sd936854, 32'sd1124278, 32'sd488820, 32'sd919949, 32'sd438893,
32'sd922215, 32'sd843131, 32'sd827901, 32'sd930301, 32'sd559519, 32'sd617543, 32'sd544751, 32'sd756909, 32'sd966568, 32'sd442012, 32'sd811494, 32'sd1085372, 32'sd787643, 32'sd958573,
32'sd958818, 32'sd774228, 32'sd857936, 32'sd625407, 32'sd963907, 32'sd854397, 32'sd1060937, 32'sd570407, 32'sd1083342, 32'sd763961, 32'sd1021194, 32'sd1164769, 32'sd448702, 32'sd1163816,
32'sd709978, 32'sd408216, 32'sd638007, 32'sd892481, 32'sd612179, 32'sd1024756, 32'sd590002, 32'sd434162, 32'sd415098, 32'sd813223, 32'sd610798, 32'sd698190, 32'sd571006, 32'sd549677,
32'sd1044186, 32'sd995487, 32'sd515913, 32'sd761323, 32'sd1206237, 32'sd874168, 32'sd736186, 32'sd708609, 32'sd791507, 32'sd677003, 32'sd856739, 32'sd686105, 32'sd516014, 32'sd618274,
32'sd1028876, 32'sd671682, 32'sd896497, 32'sd610784, 32'sd465869, 32'sd770720, 32'sd633542, 32'sd450866, 32'sd1085085, 32'sd940155, 32'sd920449, 32'sd882091, 32'sd817597, 32'sd1190557,
32'sd407624, 32'sd427795, 32'sd751877, 32'sd661599, 32'sd647016, 32'sd864661, 32'sd856419, 32'sd417758, 32'sd1105780, 32'sd624871, 32'sd1079894, 32'sd739819, 32'sd991046, 32'sd1006065,
32'sd935982, 32'sd820755, 32'sd505037, 32'sd592474, 32'sd601138, 32'sd746055, 32'sd763734, 32'sd1095767, 32'sd1038629, 32'sd503240, 32'sd478043, 32'sd731418, 32'sd898819, 32'sd508356,
32'sd1170149, 32'sd710130, 32'sd1192869, 32'sd1122039, 32'sd1196356, 32'sd436210, 32'sd693792, 32'sd1073659, 32'sd641186, 32'sd1024940, 32'sd1204657, 32'sd1158890, 32'sd1125603, 32'sd549815,
32'sd701905, 32'sd591080, 32'sd1020049, 32'sd794965, 32'sd604066, 32'sd1048641, 32'sd695558, 32'sd446360, 32'sd470421, 32'sd609912, 32'sd1201021, 32'sd887325, 32'sd816403, 32'sd1062714,
32'sd553335, 32'sd617217, 32'sd1105950, 32'sd787992, 32'sd800160, 32'sd800884, 32'sd977267, 32'sd803625, 32'sd661133, 32'sd763225, 32'sd1089736, 32'sd1175095, 32'sd714530, 32'sd977941,
32'sd539137, 32'sd532904, 32'sd981571, 32'sd598705, 32'sd448136, 32'sd532997, 32'sd890764, 32'sd1202331, 32'sd1127842, 32'sd1052209, 32'sd603071, 32'sd493962, 32'sd707028, 32'sd521575,
32'sd635902, 32'sd895239, 32'sd1189460, 32'sd576689, 32'sd731204, 32'sd939675, 32'sd467486, 32'sd977626, 32'sd842640, 32'sd866254, 32'sd594006, 32'sd883755, 32'sd1136064, 32'sd424598,
32'sd731739, 32'sd500954, 32'sd1064357, 32'sd676389, 32'sd1117396, 32'sd1171503, 32'sd791501, 32'sd646833, 32'sd620133, 32'sd795494, 32'sd762128, 32'sd1206685, 32'sd513427, 32'sd1032178,
32'sd459909, 32'sd420954, 32'sd1105954, 32'sd1125468, 32'sd1060305, 32'sd845436, 32'sd753236, 32'sd571312, 32'sd545140, 32'sd780296, 32'sd414202, 32'sd876430, 32'sd434696, 32'sd1181576,
32'sd467522, 32'sd765482, 32'sd453869, 32'sd543289, 32'sd626222, 32'sd802417, 32'sd552747, 32'sd775446, 32'sd603841, 32'sd773799, 32'sd1089263, 32'sd495497, 32'sd881257, 32'sd713811,
32'sd1171933, 32'sd422149, 32'sd974318, 32'sd1062807, 32'sd941089, 32'sd427202, 32'sd1089902, 32'sd971377, 32'sd472468, 32'sd557354, 32'sd858572, 32'sd952610, 32'sd637876, 32'sd555455,
32'sd847776, 32'sd454936, 32'sd1112818, 32'sd764743, 32'sd694729, 32'sd1022693, 32'sd579516, 32'sd586394, 32'sd484899, 32'sd664451, 32'sd631925, 32'sd884509, 32'sd928991, 32'sd951515,
32'sd1207126, 32'sd795171, 32'sd1163877, 32'sd814044, 32'sd431307, 32'sd745574, 32'sd664407, 32'sd471989, 32'sd404687, 32'sd674508, 32'sd507863, 32'sd1008217, 32'sd516180, 32'sd959980,
32'sd1089566, 32'sd843314, 32'sd605997, 32'sd988214, 32'sd682134, 32'sd514757, 32'sd885674, 32'sd1175308, 32'sd513033, 32'sd1032954, 32'sd772852, 32'sd620276, 32'sd714265, 32'sd1130482,
32'sd703834, 32'sd1192414, 32'sd987200, 32'sd568892, 32'sd713164, 32'sd528089, 32'sd1121880, 32'sd995756, 32'sd719235, 32'sd606775, 32'sd753965, 32'sd1139957, 32'sd1181692, 32'sd667069,
32'sd687699, 32'sd1078081, 32'sd1205688, 32'sd621579, 32'sd844902, 32'sd843699, 32'sd1088946, 32'sd681203, 32'sd1084952, 32'sd1144206, 32'sd761012, 32'sd581211, 32'sd918112, 32'sd467693,
32'sd819183, 32'sd1077840, 32'sd704332, 32'sd634515, 32'sd560876, 32'sd533672, 32'sd456949, 32'sd608888, 32'sd759157, 32'sd407995, 32'sd632277, 32'sd574776, 32'sd734536, 32'sd711166,
32'sd806468, 32'sd921981, 32'sd837543, 32'sd983595, 32'sd1000309, 32'sd600941, 32'sd1078841, 32'sd468510, 32'sd1085435, 32'sd431497, 32'sd942122, 32'sd877461, 32'sd511635, 32'sd457300,
32'sd935291, 32'sd770362, 32'sd909659, 32'sd593360, 32'sd578327, 32'sd797490, 32'sd999396, 32'sd585648, 32'sd684142, 32'sd1119363, 32'sd1171156, 32'sd827055, 32'sd904721, 32'sd547467,
32'sd1135843, 32'sd1042130, 32'sd692571, 32'sd441583, 32'sd701987, 32'sd608227, 32'sd1181560, 32'sd769647, 32'sd838744, 32'sd619695, 32'sd733109, 32'sd814539, 32'sd931697, 32'sd476232,
32'sd882045, 32'sd836995, 32'sd1183089, 32'sd846570, 32'sd482826, 32'sd669135, 32'sd963294, 32'sd694414, 32'sd801653, 32'sd902316, 32'sd648403, 32'sd1184482, 32'sd792531, 32'sd663271,
32'sd507927, 32'sd1072387, 32'sd431241, 32'sd655858, 32'sd1198659, 32'sd863073, 32'sd1070015, 32'sd876571, 32'sd704785, 32'sd764340, 32'sd481043, 32'sd561481, 32'sd1035612, 32'sd587211,
32'sd1047093, 32'sd999747, 32'sd490778, 32'sd787320, 32'sd456056, 32'sd678816, 32'sd403905, 32'sd826752, 32'sd735866, 32'sd636199, 32'sd519804, 32'sd1036043, 32'sd799955, 32'sd1138688,
32'sd895582, 32'sd774687, 32'sd473486, 32'sd946202, 32'sd1056966, 32'sd790299, 32'sd784506, 32'sd544689, 32'sd429684, 32'sd695103, 32'sd973732, 32'sd854959, 32'sd971383, 32'sd876747,
32'sd833860, 32'sd515302, 32'sd1041598, 32'sd430783, 32'sd433613, 32'sd1183737, 32'sd911467, 32'sd1039646, 32'sd863209, 32'sd416091, 32'sd779341, 32'sd608664, 32'sd878178, 32'sd1067941,
32'sd1137972, 32'sd745014, 32'sd1041245, 32'sd971802, 32'sd642511, 32'sd626436, 32'sd887915, 32'sd913796, 32'sd572181, 32'sd1106988, 32'sd1194625, 32'sd548421, 32'sd880955, 32'sd747452,
32'sd1167861, 32'sd417065, 32'sd1069394, 32'sd526384, 32'sd716362, 32'sd662331, 32'sd1073043, 32'sd854287, 32'sd827478, 32'sd1009588, 32'sd884706, 32'sd545751, 32'sd974402, 32'sd663644,
32'sd1052348, 32'sd699955, 32'sd805481, 32'sd1106045, 32'sd1068407, 32'sd842160, 32'sd1018699, 32'sd827863, 32'sd897148, 32'sd594229, 32'sd1115336, 32'sd747056, 32'sd1052035, 32'sd407625,
32'sd855644, 32'sd795536, 32'sd458469, 32'sd536513, 32'sd746757, 32'sd958933, 32'sd442522, 32'sd513321, 32'sd998883, 32'sd776422, 32'sd906731, 32'sd1017555, 32'sd1132635, 32'sd621089,
32'sd910252, 32'sd1110147, 32'sd1129418, 32'sd870058, 32'sd797410, 32'sd1032997, 32'sd1108323, 32'sd1189962, 32'sd1172786, 32'sd507964, 32'sd598368, 32'sd429735, 32'sd1119782, 32'sd864056,
32'sd985506, 32'sd1078719, 32'sd692547, 32'sd937396, 32'sd784267, 32'sd1046097, 32'sd691583, 32'sd1168631, 32'sd545769, 32'sd509257, 32'sd561392, 32'sd1126145, 32'sd702470, 32'sd1051780,
32'sd680771, 32'sd767912, 32'sd842576, 32'sd1205813, 32'sd427390, 32'sd786258, 32'sd503730, 32'sd961618, 32'sd661497, 32'sd1176025, 32'sd852393, 32'sd664262, 32'sd875439, 32'sd1132651,
32'sd1131713, 32'sd1000923, 32'sd997553, 32'sd576987, 32'sd519213, 32'sd668903, 32'sd433379, 32'sd695203, 32'sd884181, 32'sd1130633, 32'sd653238, 32'sd522616, 32'sd968701, 32'sd1145731,
32'sd757250, 32'sd918858, 32'sd1118882, 32'sd685904, 32'sd1142963, 32'sd663430, 32'sd432158, 32'sd1134148, 32'sd1178480, 32'sd562958, 32'sd1010202, 32'sd429702, 32'sd1204621, 32'sd520576,
32'sd719728, 32'sd415784, 32'sd523064, 32'sd1091282, 32'sd660358, 32'sd510520, 32'sd911756, 32'sd496082, 32'sd723046, 32'sd1145917, 32'sd823646, 32'sd1057909, 32'sd902613, 32'sd593769,
32'sd895952, 32'sd896462, 32'sd1051056, 32'sd437478, 32'sd965386, 32'sd917870, 32'sd469068, 32'sd669213, 32'sd894242, 32'sd466288, 32'sd990888, 32'sd981434, 32'sd554534, 32'sd855929,
32'sd1162652, 32'sd761132, 32'sd1117118, 32'sd677971, 32'sd1201164, 32'sd1076968, 32'sd622828, 32'sd1119081, 32'sd660204, 32'sd880177, 32'sd560847, 32'sd919405, 32'sd566525, 32'sd1068826,
32'sd795601, 32'sd691463, 32'sd842009, 32'sd581274, 32'sd685141, 32'sd671852, 32'sd1039824, 32'sd681553, 32'sd611952, 32'sd1054833, 32'sd790448, 32'sd989629, 32'sd995366, 32'sd976315,
32'sd1153129, 32'sd650095, 32'sd793560, 32'sd491928, 32'sd1053598, 32'sd678470, 32'sd632149, 32'sd479190, 32'sd642780, 32'sd432024, 32'sd778379, 32'sd1047702, 32'sd553321, 32'sd847715,
32'sd891940, 32'sd574860, 32'sd625846, 32'sd754919, 32'sd920466, 32'sd790495, 32'sd1160846, 32'sd859296, 32'sd512105, 32'sd925851, 32'sd669871, 32'sd1061438, 32'sd524590, 32'sd1152554,
32'sd619233, 32'sd956536, 32'sd912122, 32'sd846903, 32'sd1129105, 32'sd1193145, 32'sd883141, 32'sd768700, 32'sd983251, 32'sd1158901, 32'sd915666, 32'sd676180, 32'sd712538, 32'sd1181316,
32'sd476558, 32'sd1101430, 32'sd585147, 32'sd427362, 32'sd771959, 32'sd571146, 32'sd1072861, 32'sd496873, 32'sd620237, 32'sd1125813, 32'sd699471, 32'sd796284, 32'sd1047886, 32'sd928028,
32'sd772168, 32'sd619602, 32'sd592116, 32'sd1163659, 32'sd599796, 32'sd494592, 32'sd549489, 32'sd1024312, 32'sd730219, 32'sd1096551, 32'sd1110638, 32'sd567179, 32'sd996964, 32'sd1012185,
32'sd729554, 32'sd1100880, 32'sd792314, 32'sd532948, 32'sd642573, 32'sd901739, 32'sd482208, 32'sd414713, 32'sd757002, 32'sd1156524, 32'sd582492, 32'sd463723, 32'sd408702, 32'sd954764,
32'sd590246, 32'sd1207084, 32'sd803109, 32'sd453735, 32'sd904651, 32'sd926048, 32'sd1119478, 32'sd938332, 32'sd654990, 32'sd953943, 32'sd870999, 32'sd1086760, 32'sd921069, 32'sd782067,
32'sd649486, 32'sd696438, 32'sd812770, 32'sd792845, 32'sd693759, 32'sd648449, 32'sd1140466, 32'sd935577, 32'sd899745, 32'sd956613, 32'sd1162861, 32'sd1119362, 32'sd984541, 32'sd659714,
32'sd1033733, 32'sd608539, 32'sd443805, 32'sd923278, 32'sd989868, 32'sd1154663, 32'sd405928, 32'sd893874, 32'sd1053737, 32'sd595207, 32'sd1189910, 32'sd582188, 32'sd1139332, 32'sd794561,
32'sd597681, 32'sd432055, 32'sd1068426, 32'sd919199, 32'sd492175, 32'sd933504, 32'sd1037852, 32'sd741106, 32'sd834121, 32'sd594947, 32'sd589792, 32'sd1018947, 32'sd952123, 32'sd824966,
32'sd539967, 32'sd508694, 32'sd694030, 32'sd745578, 32'sd1105929, 32'sd929267, 32'sd1049238, 32'sd671948, 32'sd1132043, 32'sd648785, 32'sd984693, 32'sd1186579, 32'sd1177248, 32'sd720882,
32'sd542733, 32'sd1109640, 32'sd1073414, 32'sd608409, 32'sd568956, 32'sd899292, 32'sd641110, 32'sd686232, 32'sd1197025, 32'sd632108, 32'sd1155632, 32'sd786679, 32'sd957435, 32'sd501087,
32'sd533788, 32'sd1108622, 32'sd963656, 32'sd447702, 32'sd739033, 32'sd407537, 32'sd856750, 32'sd528861, 32'sd587827, 32'sd592741, 32'sd947438, 32'sd993578, 32'sd540985, 32'sd627754,
32'sd597399, 32'sd1207951, 32'sd424448, 32'sd702085, 32'sd886813, 32'sd555862, 32'sd706021, 32'sd672985, 32'sd1101978, 32'sd1167927, 32'sd734590, 32'sd409897, 32'sd1166738, 32'sd571776,
32'sd1208094, 32'sd841286, 32'sd526705, 32'sd729540, 32'sd1115131, 32'sd505240, 32'sd867607, 32'sd735250, 32'sd581486, 32'sd488365, 32'sd686268, 32'sd984363, 32'sd937910, 32'sd1140173,
32'sd798033, 32'sd1150440, 32'sd764558, 32'sd427174, 32'sd761324, 32'sd928750, 32'sd1028768, 32'sd1141269, 32'sd539287, 32'sd688630, 32'sd764858, 32'sd1139365, 32'sd841411, 32'sd915020,
32'sd525850, 32'sd679644, 32'sd1057495, 32'sd773351, 32'sd574715, 32'sd905551, 32'sd549755, 32'sd576508, 32'sd685507, 32'sd707883, 32'sd1093163, 32'sd492046, 32'sd1101877, 32'sd951089,
32'sd1092191, 32'sd921183, 32'sd873019, 32'sd1074512, 32'sd526559, 32'sd1040818, 32'sd1073818, 32'sd474116, 32'sd667808, 32'sd1201235, 32'sd802850, 32'sd989301, 32'sd423385, 32'sd463549,
32'sd782197, 32'sd815536, 32'sd1175160, 32'sd1082582, 32'sd966812, 32'sd960157, 32'sd1018621, 32'sd889775, 32'sd1196951, 32'sd478047, 32'sd746383, 32'sd448743, 32'sd943333, 32'sd1065750,
32'sd985437, 32'sd856032, 32'sd637904, 32'sd1069014, 32'sd527013, 32'sd798587, 32'sd442618, 32'sd1198654, 32'sd541720, 32'sd960291, 32'sd527105, 32'sd444731, 32'sd539236, 32'sd535723,
32'sd896930, 32'sd577085, 32'sd617545, 32'sd649555, 32'sd815290, 32'sd927906, 32'sd902593, 32'sd858930, 32'sd864605, 32'sd1108817, 32'sd845531, 32'sd873249, 32'sd629543, 32'sd618567,
32'sd646820, 32'sd781646, 32'sd816485, 32'sd642903, 32'sd672302, 32'sd793930, 32'sd605520, 32'sd968757, 32'sd690309, 32'sd1071707, 32'sd545848, 32'sd643089, 32'sd1174112, 32'sd1183484,
32'sd747644, 32'sd617299, 32'sd1207592, 32'sd984795, 32'sd987273, 32'sd1017541, 32'sd606043, 32'sd1141637, 32'sd430034, 32'sd900951, 32'sd1209165, 32'sd951347, 32'sd880887, 32'sd512788,
32'sd456931, 32'sd949652, 32'sd632962, 32'sd640090, 32'sd582490, 32'sd1136194, 32'sd686305, 32'sd1206106, 32'sd737384, 32'sd861777, 32'sd1153146, 32'sd546034, 32'sd586792, 32'sd852889,
32'sd509823, 32'sd456117, 32'sd488862, 32'sd854938, 32'sd1186455, 32'sd785801, 32'sd1007768, 32'sd650380, 32'sd732754, 32'sd621460, 32'sd726870, 32'sd918238, 32'sd851489, 32'sd1072771,
32'sd792026, 32'sd520858, 32'sd819947, 32'sd1012892, 32'sd1078785, 32'sd1124723, 32'sd974163, 32'sd680582, 32'sd732072, 32'sd1016111, 32'sd723714, 32'sd707960, 32'sd834557, 32'sd546106,
32'sd856345, 32'sd630408, 32'sd586628, 32'sd721689, 32'sd995550, 32'sd737949, 32'sd1118191, 32'sd865892, 32'sd773862, 32'sd583371, 32'sd551402, 32'sd986491, 32'sd764262, 32'sd842824,
32'sd745668, 32'sd1128642, 32'sd804600, 32'sd655480, 32'sd931359, 32'sd927316, 32'sd855270, 32'sd824379, 32'sd780354, 32'sd1104870, 32'sd1142395, 32'sd1018608, 32'sd766497, 32'sd719361,
32'sd856237, 32'sd559063, 32'sd1011056, 32'sd919857, 32'sd1120962, 32'sd800723, 32'sd799920, 32'sd493498, 32'sd1016362, 32'sd469793, 32'sd1104438, 32'sd558986, 32'sd1090793, 32'sd1207793,
32'sd665382, 32'sd473530, 32'sd887034, 32'sd1004847, 32'sd512847, 32'sd885350, 32'sd597303, 32'sd857055, 32'sd1041661, 32'sd1046491, 32'sd452328, 32'sd924789, 32'sd1007764, 32'sd1038873,
32'sd1015577, 32'sd878388, 32'sd663542, 32'sd411206, 32'sd885811, 32'sd467221, 32'sd444333, 32'sd672897, 32'sd1024502, 32'sd724930, 32'sd858962, 32'sd642332, 32'sd995223, 32'sd798863,
32'sd1182067, 32'sd905861, 32'sd563196, 32'sd540078, 32'sd516678, 32'sd821805, 32'sd844300, 32'sd464132, 32'sd970516, 32'sd1115947, 32'sd1150514, 32'sd625226, 32'sd1028372, 32'sd534493,
32'sd493193, 32'sd413372, 32'sd951475, 32'sd615260, 32'sd920023, 32'sd769998, 32'sd745465, 32'sd1194860, 32'sd1160956, 32'sd1179848, 32'sd821729, 32'sd999236, 32'sd1073938, 32'sd754947,
32'sd460315, 32'sd636493, 32'sd1175642, 32'sd1127679, 32'sd843753, 32'sd1034034, 32'sd1187407, 32'sd1152415, 32'sd413467, 32'sd787742, 32'sd964779, 32'sd1078948, 32'sd572482, 32'sd552323,
32'sd1015784, 32'sd665584, 32'sd1104055, 32'sd765740, 32'sd779658, 32'sd504799, 32'sd514088, 32'sd743545, 32'sd836900, 32'sd1082384, 32'sd821088, 32'sd888819, 32'sd568679, 32'sd1047018,
32'sd935181, 32'sd1165600, 32'sd684467, 32'sd932993, 32'sd1178646, 32'sd814387, 32'sd884457, 32'sd1021944, 32'sd998678, 32'sd1208933, 32'sd837160, 32'sd1004510, 32'sd1077548, 32'sd763157,
32'sd627726, 32'sd742849, 32'sd913458, 32'sd800162, 32'sd514840, 32'sd1085434, 32'sd961327, 32'sd553884, 32'sd894971, 32'sd784231, 32'sd867655, 32'sd598991, 32'sd1028409, 32'sd1139842,
32'sd1154562, 32'sd1139631, 32'sd710240, 32'sd645364, 32'sd900088, 32'sd496129, 32'sd568534, 32'sd1101404, 32'sd1143623, 32'sd956627, 32'sd923491, 32'sd710787, 32'sd720636, 32'sd1106124,
32'sd853102, 32'sd957772, 32'sd876222, 32'sd888269, 32'sd1178072, 32'sd463900, 32'sd1136666, 32'sd569286, 32'sd687651, 32'sd1070547, 32'sd604040, 32'sd629628, 32'sd519886, 32'sd1187854,
32'sd962743, 32'sd883273, 32'sd416523, 32'sd576916, 32'sd849518, 32'sd927666, 32'sd1049747, 32'sd901658, 32'sd1131695, 32'sd892032, 32'sd1191139, 32'sd607038, 32'sd1081810, 32'sd1179903,
32'sd725055, 32'sd1166077, 32'sd761153, 32'sd561571, 32'sd519022, 32'sd1148425, 32'sd728986, 32'sd890231, 32'sd639102, 32'sd752893, 32'sd1189271, 32'sd891151, 32'sd1165454, 32'sd999813,
32'sd738335, 32'sd650180, 32'sd935543, 32'sd1017511, 32'sd496887, 32'sd422828, 32'sd991885, 32'sd424247, 32'sd661448, 32'sd702865, 32'sd1025302, 32'sd446308, 32'sd1104183, 32'sd814093,
32'sd1197367, 32'sd874607, 32'sd981751, 32'sd953022, 32'sd406607, 32'sd720181, 32'sd1196223, 32'sd534781, 32'sd722233, 32'sd586077, 32'sd1169048, 32'sd1101989, 32'sd1167736, 32'sd566538,
32'sd692297, 32'sd710497, 32'sd479562, 32'sd504727, 32'sd1178067, 32'sd1108436, 32'sd968439, 32'sd1127894, 32'sd635118, 32'sd588058, 32'sd710734, 32'sd453474, 32'sd1079928, 32'sd821980,
32'sd918482, 32'sd656035, 32'sd939085, 32'sd1184963, 32'sd690467, 32'sd1113576, 32'sd891468, 32'sd673351, 32'sd950648, 32'sd894291, 32'sd624306, 32'sd596995, 32'sd1130710, 32'sd1208402,
32'sd1053114, 32'sd420724, 32'sd1157599, 32'sd550281, 32'sd584720, 32'sd1070469, 32'sd468274, 32'sd824383, 32'sd598712, 32'sd690766, 32'sd1197843, 32'sd479630, 32'sd930310, 32'sd1131654,
32'sd912225, 32'sd905422, 32'sd462516, 32'sd703856, 32'sd706042, 32'sd925118, 32'sd878378, 32'sd938755, 32'sd1197500, 32'sd670077, 32'sd923247, 32'sd1146265, 32'sd956277, 32'sd1015870,
32'sd659158, 32'sd856785, 32'sd789815, 32'sd671378, 32'sd511371, 32'sd968380, 32'sd1012902, 32'sd717992, 32'sd693382, 32'sd1039301, 32'sd1000965, 32'sd855947, 32'sd987541, 32'sd741984,
32'sd443419, 32'sd1038066, 32'sd824799, 32'sd708521, 32'sd799297, 32'sd1127639, 32'sd1003954, 32'sd717066, 32'sd538385, 32'sd908005, 32'sd924632, 32'sd990599, 32'sd509235, 32'sd755395,
32'sd755971, 32'sd918911, 32'sd857035, 32'sd564889, 32'sd918633, 32'sd1170841, 32'sd633404, 32'sd431306, 32'sd754801, 32'sd983208, 32'sd624657, 32'sd657780, 32'sd671450, 32'sd523069,
32'sd878124, 32'sd1071080, 32'sd1083580, 32'sd1048430, 32'sd689132, 32'sd409713, 32'sd1085457, 32'sd1091814, 32'sd893299, 32'sd915393, 32'sd1201863, 32'sd728207, 32'sd1030659, 32'sd817273,
32'sd1171523, 32'sd1183573, 32'sd559667, 32'sd1016162, 32'sd564861, 32'sd658150, 32'sd484806, 32'sd681909, 32'sd442477, 32'sd924695, 32'sd441636, 32'sd826140, 32'sd1026057, 32'sd595790,
32'sd969088, 32'sd976771, 32'sd1180799, 32'sd718486, 32'sd1207022, 32'sd757995, 32'sd1208301, 32'sd598579, 32'sd735175, 32'sd613165, 32'sd471887, 32'sd450088, 32'sd635863, 32'sd922710,
32'sd909247, 32'sd545203, 32'sd1204260, 32'sd701056, 32'sd1023295, 32'sd416819, 32'sd508882, 32'sd1130818, 32'sd744876, 32'sd1037990, 32'sd1182669, 32'sd819665, 32'sd1079589, 32'sd771239,
32'sd865372, 32'sd637635, 32'sd977789, 32'sd1127554, 32'sd507536, 32'sd698456, 32'sd796982, 32'sd997598, 32'sd1133710, 32'sd748811, 32'sd1087103, 32'sd454252, 32'sd660886, 32'sd664325,
32'sd690166, 32'sd587463, 32'sd414450, 32'sd690368, 32'sd505278, 32'sd927292, 32'sd570714, 32'sd770843, 32'sd632595, 32'sd1034888, 32'sd938924, 32'sd614660, 32'sd975490, 32'sd440870,
32'sd1006943, 32'sd1097729, 32'sd536069, 32'sd1190675, 32'sd683297, 32'sd852768, 32'sd493824, 32'sd465223, 32'sd405516, 32'sd598517, 32'sd405352, 32'sd453262, 32'sd604189, 32'sd765470,
32'sd529535, 32'sd1015767, 32'sd585759, 32'sd805699, 32'sd750443, 32'sd794953, 32'sd577869, 32'sd1052905, 32'sd1120603, 32'sd845163, 32'sd411730, 32'sd643576, 32'sd1042001, 32'sd698799,
32'sd404811, 32'sd699245, 32'sd546238, 32'sd886526, 32'sd446373, 32'sd745229, 32'sd859056, 32'sd1009437, 32'sd946326, 32'sd800417, 32'sd1193744, 32'sd950867, 32'sd933873, 32'sd502199,
32'sd436143, 32'sd970065, 32'sd582501, 32'sd1202849, 32'sd569232, 32'sd800316, 32'sd1068850, 32'sd1031939, 32'sd612868, 32'sd557222, 32'sd795922, 32'sd893610, 32'sd748490, 32'sd951945,
32'sd596605, 32'sd712863, 32'sd1075356, 32'sd565433, 32'sd966521, 32'sd1174895, 32'sd704050, 32'sd527759, 32'sd889346, 32'sd750873, 32'sd545213, 32'sd547741, 32'sd1045390, 32'sd591274,
32'sd801373, 32'sd842713, 32'sd1167483, 32'sd404995, 32'sd439923, 32'sd787983, 32'sd807551, 32'sd1004475, 32'sd405841, 32'sd1165790, 32'sd1021743, 32'sd926381, 32'sd512353, 32'sd431836,
32'sd864536, 32'sd1088606, 32'sd629594, 32'sd1159685, 32'sd1004159, 32'sd488134, 32'sd476457, 32'sd1164056, 32'sd900523, 32'sd1117051, 32'sd1040136, 32'sd638431, 32'sd1100121, 32'sd472248,
32'sd1175485, 32'sd574143, 32'sd680980, 32'sd769419, 32'sd519297, 32'sd875019, 32'sd885565, 32'sd438248, 32'sd924371, 32'sd1177320, 32'sd685744, 32'sd1121832, 32'sd570165, 32'sd1018126,
32'sd753637, 32'sd644399, 32'sd613831, 32'sd925648, 32'sd435050, 32'sd1063451, 32'sd639404, 32'sd588259, 32'sd517144, 32'sd1065722, 32'sd826580, 32'sd701155, 32'sd830230, 32'sd433653,
32'sd661379, 32'sd528589, 32'sd771960, 32'sd866805, 32'sd478431, 32'sd633547, 32'sd1178306, 32'sd1183624, 32'sd788161, 32'sd716113, 32'sd930488, 32'sd493874, 32'sd900052, 32'sd1123118,
32'sd446875, 32'sd767088, 32'sd825963, 32'sd491071, 32'sd1100029, 32'sd931031, 32'sd564817, 32'sd505346, 32'sd960390, 32'sd809474, 32'sd1051383, 32'sd858408, 32'sd899329, 32'sd821366,
32'sd796854, 32'sd898134, 32'sd695445, 32'sd861761, 32'sd518114, 32'sd502618, 32'sd609256, 32'sd457095, 32'sd696984, 32'sd741303, 32'sd723778, 32'sd835508, 32'sd580456, 32'sd1115080,
32'sd1191939, 32'sd797234, 32'sd1034965, 32'sd1048491, 32'sd1115268, 32'sd916159, 32'sd898985, 32'sd990497, 32'sd464367, 32'sd573723, 32'sd1126832, 32'sd1072008, 32'sd618066, 32'sd902930,
32'sd1022996, 32'sd781931, 32'sd930591, 32'sd632637, 32'sd452453, 32'sd1190867, 32'sd1198861, 32'sd504224, 32'sd855760, 32'sd838157, 32'sd1096986, 32'sd994804, 32'sd1158783, 32'sd975476,
32'sd844479, 32'sd970630, 32'sd690813, 32'sd737204, 32'sd497342, 32'sd955302, 32'sd939940, 32'sd1110174, 32'sd496269, 32'sd574601, 32'sd537562, 32'sd475418, 32'sd940040, 32'sd719755,
32'sd990875, 32'sd663262, 32'sd1094935, 32'sd832527, 32'sd1053494, 32'sd976973, 32'sd756517, 32'sd543997, 32'sd1143158, 32'sd1077238, 32'sd795151, 32'sd865377, 32'sd652782, 32'sd526511,
32'sd791364, 32'sd646208, 32'sd963259, 32'sd947608, 32'sd932861, 32'sd663133, 32'sd437383, 32'sd530520, 32'sd616634, 32'sd1089895, 32'sd1083066, 32'sd990878, 32'sd1175392, 32'sd1121852,
32'sd1054650, 32'sd882576, 32'sd1134422, 32'sd1095031, 32'sd485408, 32'sd1066495, 32'sd1162366, 32'sd612255, 32'sd568936, 32'sd964438, 32'sd841996, 32'sd628320, 32'sd823326, 32'sd428962,
32'sd555439, 32'sd662268, 32'sd755520, 32'sd548516, 32'sd594445, 32'sd524060, 32'sd920054, 32'sd636720, 32'sd808000, 32'sd661339, 32'sd606440, 32'sd405332, 32'sd838252, 32'sd1177566,
32'sd993617, 32'sd861071, 32'sd645793, 32'sd460573, 32'sd520715, 32'sd1123324, 32'sd463856, 32'sd960975, 32'sd505241, 32'sd712727, 32'sd962343, 32'sd688898, 32'sd455211, 32'sd520023,
32'sd997662, 32'sd713333, 32'sd854326, 32'sd1092292, 32'sd687827, 32'sd473677, 32'sd653954, 32'sd1205529, 32'sd1010405, 32'sd1056553, 32'sd656234, 32'sd597997, 32'sd761314, 32'sd563256,
32'sd622936, 32'sd1084904, 32'sd983289, 32'sd579244, 32'sd557374, 32'sd755417, 32'sd1197833, 32'sd600528, 32'sd1172698, 32'sd1204145, 32'sd962690, 32'sd1107525, 32'sd1063706, 32'sd874037,
32'sd534815, 32'sd713497, 32'sd888741, 32'sd1133370, 32'sd1047567, 32'sd750550, 32'sd806323, 32'sd447839, 32'sd985488, 32'sd562367, 32'sd1073711, 32'sd674086, 32'sd784017, 32'sd1109430,
32'sd623883, 32'sd542911, 32'sd663672, 32'sd1154889, 32'sd1083878, 32'sd764193, 32'sd1046150, 32'sd892008, 32'sd740387, 32'sd848520, 32'sd489491, 32'sd752218, 32'sd697710, 32'sd1011369,
32'sd773333, 32'sd500116, 32'sd887377, 32'sd453367, 32'sd554811, 32'sd1148927, 32'sd655448, 32'sd1161775, 32'sd523894, 32'sd822609, 32'sd845136, 32'sd775461, 32'sd673936, 32'sd1138259,
32'sd834475, 32'sd598952, 32'sd1177573, 32'sd834315, 32'sd673212, 32'sd637726, 32'sd1193925, 32'sd804591, 32'sd1053869, 32'sd1154641, 32'sd1172645, 32'sd426915, 32'sd918489, 32'sd455772,
32'sd1106625, 32'sd527507, 32'sd1031081, 32'sd766203, 32'sd1143126, 32'sd578353, 32'sd1096485, 32'sd1149973, 32'sd1048576, 32'sd627029, 32'sd1003774, 32'sd586351, 32'sd895325, 32'sd822739,
32'sd859723, 32'sd1188735, 32'sd571650, 32'sd790063, 32'sd737605, 32'sd666858, 32'sd714988, 32'sd1040316, 32'sd458849, 32'sd648681, 32'sd699449, 32'sd706856, 32'sd914913, 32'sd857272,
32'sd973751, 32'sd1014886, 32'sd1183837, 32'sd817098, 32'sd1047778, 32'sd866217, 32'sd817387, 32'sd1100448, 32'sd779205, 32'sd426866, 32'sd795871, 32'sd503334, 32'sd509127, 32'sd486983,
32'sd466782, 32'sd683546, 32'sd853456, 32'sd517379, 32'sd867345, 32'sd795880, 32'sd886693, 32'sd939969, 32'sd922592, 32'sd439674, 32'sd1055374, 32'sd1091715, 32'sd972098, 32'sd1102061,
32'sd977226, 32'sd1154160, 32'sd973737, 32'sd721866, 32'sd508620, 32'sd1032524, 32'sd1018190, 32'sd856723, 32'sd495500, 32'sd1140503, 32'sd973955, 32'sd1207201, 32'sd530149, 32'sd427387,
32'sd1044244, 32'sd893735, 32'sd655105, 32'sd984322, 32'sd1038253, 32'sd1101491, 32'sd864888, 32'sd1144622, 32'sd1090151, 32'sd1079372, 32'sd453656, 32'sd802490, 32'sd900353, 32'sd836440,
32'sd645735, 32'sd821116, 32'sd1193503, 32'sd585472, 32'sd1108346, 32'sd641414, 32'sd472272, 32'sd772915, 32'sd891603, 32'sd538350, 32'sd522161, 32'sd1061566, 32'sd906946, 32'sd582615,
32'sd873091, 32'sd800607, 32'sd564055, 32'sd859166, 32'sd1066478, 32'sd804619, 32'sd823191, 32'sd1074568, 32'sd755292, 32'sd433732, 32'sd873442, 32'sd523739, 32'sd919735, 32'sd1192148,
32'sd1107786, 32'sd529576, 32'sd453360, 32'sd844653, 32'sd706405, 32'sd749191, 32'sd1056304, 32'sd1021649, 32'sd1187402, 32'sd1183940, 32'sd1164618, 32'sd542618, 32'sd832660, 32'sd462201,
32'sd636569, 32'sd573269, 32'sd847448, 32'sd403777, 32'sd458101, 32'sd861289, 32'sd708048, 32'sd770171, 32'sd630276, 32'sd1136441, 32'sd739823, 32'sd1124653, 32'sd1093893, 32'sd991750,
32'sd572729, 32'sd734323, 32'sd815222, 32'sd1103276, 32'sd934179, 32'sd814893, 32'sd636064, 32'sd1178509, 32'sd415951, 32'sd909809, 32'sd669582, 32'sd674104, 32'sd586606, 32'sd660637,
32'sd1137302, 32'sd715279, 32'sd759195, 32'sd429529, 32'sd1205017, 32'sd1023956, 32'sd1087520, 32'sd683464, 32'sd1075024, 32'sd820967, 32'sd692654, 32'sd770586, 32'sd1043605, 32'sd777099,
32'sd1024113, 32'sd765167, 32'sd506651, 32'sd451220, 32'sd545556, 32'sd973159, 32'sd578167, 32'sd996030, 32'sd994783, 32'sd1152199, 32'sd1185169, 32'sd893072, 32'sd619540, 32'sd715718,
32'sd921385, 32'sd676840, 32'sd716871, 32'sd626077, 32'sd473978, 32'sd930140, 32'sd681898, 32'sd896418, 32'sd468057, 32'sd841112, 32'sd616628, 32'sd1136012, 32'sd713818, 32'sd1130421,
32'sd565615, 32'sd1032305, 32'sd1073537, 32'sd1017097, 32'sd823365, 32'sd1161065, 32'sd845128, 32'sd569870, 32'sd1167315, 32'sd826870, 32'sd934729, 32'sd911639, 32'sd769450, 32'sd923996,
32'sd1096394, 32'sd904091, 32'sd1055534, 32'sd782932, 32'sd962779, 32'sd687839, 32'sd791695, 32'sd446074, 32'sd761302, 32'sd809140, 32'sd801135, 32'sd836464, 32'sd987567, 32'sd776962,
32'sd809396, 32'sd833269, 32'sd723228, 32'sd1185358, 32'sd795265, 32'sd997386, 32'sd1092023, 32'sd966457, 32'sd755570, 32'sd1157306, 32'sd479928, 32'sd979238, 32'sd1186305, 32'sd682318,
32'sd439230, 32'sd659198, 32'sd449599, 32'sd415009, 32'sd499575, 32'sd1064160, 32'sd901984, 32'sd765177, 32'sd477286, 32'sd891929, 32'sd1002189, 32'sd1121800, 32'sd465002, 32'sd424469,
32'sd446290, 32'sd593396, 32'sd1153307, 32'sd1059532, 32'sd693050, 32'sd1057673, 32'sd934217, 32'sd493512, 32'sd587538, 32'sd404932, 32'sd763740, 32'sd968394, 32'sd1012363, 32'sd515393,
32'sd650286, 32'sd808171, 32'sd562601, 32'sd673324, 32'sd580736, 32'sd1206705, 32'sd1172419, 32'sd602155, 32'sd1048594, 32'sd597767, 32'sd734660, 32'sd824942, 32'sd430970, 32'sd739664,
32'sd722663, 32'sd1063749, 32'sd1031801, 32'sd548309, 32'sd697419, 32'sd811355, 32'sd1108882, 32'sd712275, 32'sd984611, 32'sd692542, 32'sd471321, 32'sd538074, 32'sd656259, 32'sd426808,
32'sd1174502, 32'sd638708, 32'sd1011837, 32'sd910028, 32'sd808859, 32'sd638705, 32'sd1049674, 32'sd843205, 32'sd845448, 32'sd792338, 32'sd546064, 32'sd928710, 32'sd459461, 32'sd1151714,
32'sd461668, 32'sd549368, 32'sd1133585, 32'sd533110, 32'sd782953, 32'sd1011601, 32'sd1190095, 32'sd715669, 32'sd828248, 32'sd1138762, 32'sd418875, 32'sd541661, 32'sd1209301, 32'sd1051409,
32'sd958224, 32'sd1183478, 32'sd1112365, 32'sd947832, 32'sd775629, 32'sd1018291, 32'sd858482, 32'sd492039, 32'sd1183937, 32'sd1080309, 32'sd818056, 32'sd1038085, 32'sd831423, 32'sd947058,
32'sd848422, 32'sd1096261, 32'sd1152098, 32'sd1029020, 32'sd1118134, 32'sd678258, 32'sd1008447, 32'sd682203, 32'sd948638, 32'sd1097523, 32'sd611140, 32'sd612035, 32'sd425648, 32'sd969655,
32'sd1014222, 32'sd478502, 32'sd452196, 32'sd886886, 32'sd628783, 32'sd665588, 32'sd414735, 32'sd1068651, 32'sd957099, 32'sd481957, 32'sd516993, 32'sd470304, 32'sd837771, 32'sd1123365,
32'sd414031, 32'sd635283, 32'sd1157271, 32'sd599785, 32'sd509356, 32'sd961885, 32'sd1170764, 32'sd606785, 32'sd457301, 32'sd645351, 32'sd678428, 32'sd1048236, 32'sd742495, 32'sd666513,
32'sd1055981, 32'sd999600, 32'sd921168, 32'sd410832, 32'sd651595, 32'sd938149, 32'sd1053150, 32'sd788363, 32'sd687050, 32'sd491727, 32'sd986180, 32'sd1069452, 32'sd1151988, 32'sd1047323,
32'sd643084, 32'sd640593, 32'sd987690, 32'sd783793, 32'sd983466, 32'sd926592, 32'sd835372, 32'sd535427, 32'sd788392, 32'sd723326, 32'sd939347, 32'sd1018603, 32'sd910785, 32'sd926381,
32'sd774721, 32'sd863815, 32'sd839308, 32'sd430212, 32'sd826588, 32'sd1075601, 32'sd910904, 32'sd962330, 32'sd695427, 32'sd817523, 32'sd1116383, 32'sd693322, 32'sd706777, 32'sd536646,
32'sd554079, 32'sd1168422, 32'sd710227, 32'sd444651, 32'sd901529, 32'sd957005, 32'sd539059, 32'sd654319, 32'sd421743, 32'sd1093687, 32'sd1038447, 32'sd902951, 32'sd809299, 32'sd512953,
32'sd559687, 32'sd1118788, 32'sd795623, 32'sd439211, 32'sd835311, 32'sd868059, 32'sd873842, 32'sd926535, 32'sd1163408, 32'sd1026487, 32'sd1025589, 32'sd1025216, 32'sd661249, 32'sd1182145,
32'sd1179077, 32'sd1096053, 32'sd491618, 32'sd1139223, 32'sd821981, 32'sd1190558, 32'sd897594, 32'sd1017095, 32'sd773322, 32'sd895622, 32'sd1106396, 32'sd601670, 32'sd1005208, 32'sd622165,
32'sd418656, 32'sd572676, 32'sd668190, 32'sd990073, 32'sd812527, 32'sd451684, 32'sd1100076, 32'sd745617, 32'sd990414, 32'sd729384, 32'sd1078421, 32'sd462051, 32'sd551219, 32'sd472609,
32'sd740923, 32'sd966553, 32'sd1022549, 32'sd517381, 32'sd790382, 32'sd1097113, 32'sd1203318, 32'sd566951, 32'sd463458, 32'sd823326, 32'sd774410, 32'sd731306, 32'sd523754, 32'sd677878,
32'sd1000371, 32'sd977733, 32'sd526481, 32'sd1131932, 32'sd649059, 32'sd977026, 32'sd951691, 32'sd833605, 32'sd695193, 32'sd674513, 32'sd626264, 32'sd470905, 32'sd1077678, 32'sd1077445,
32'sd999292, 32'sd1001341, 32'sd964631, 32'sd1074520, 32'sd641203, 32'sd1123464, 32'sd807667, 32'sd758462, 32'sd618562, 32'sd706491, 32'sd454289, 32'sd1149437, 32'sd962341, 32'sd1013621,
32'sd434078, 32'sd781965, 32'sd791082, 32'sd879690, 32'sd865596, 32'sd460158, 32'sd1037198, 32'sd906247, 32'sd1017734, 32'sd463112, 32'sd625534, 32'sd730285, 32'sd763397, 32'sd942280,
32'sd1024446, 32'sd864237, 32'sd1090390, 32'sd819751, 32'sd609281, 32'sd1065395, 32'sd1122545, 32'sd609987, 32'sd635089, 32'sd689302, 32'sd1103753, 32'sd1181959, 32'sd873246, 32'sd454496,
32'sd653349, 32'sd1021857, 32'sd688832, 32'sd519543, 32'sd580423, 32'sd826886, 32'sd637669, 32'sd1186776, 32'sd823837, 32'sd926752, 32'sd486688, 32'sd626116, 32'sd897077, 32'sd1156723,
32'sd477223, 32'sd765976, 32'sd1169850, 32'sd987759, 32'sd1184905, 32'sd975926, 32'sd706739, 32'sd1010890, 32'sd910456, 32'sd1181008, 32'sd900498, 32'sd909645, 32'sd990353, 32'sd1026648,
32'sd1046324, 32'sd612789, 32'sd1142018, 32'sd423664, 32'sd868453, 32'sd1113462, 32'sd853427, 32'sd439294, 32'sd783492, 32'sd1126628, 32'sd502774, 32'sd485072, 32'sd986667, 32'sd1074569,
32'sd935463, 32'sd704134, 32'sd816075, 32'sd1012246, 32'sd599491, 32'sd1031762, 32'sd1019320, 32'sd1024132, 32'sd417228, 32'sd872844, 32'sd996041, 32'sd1132975, 32'sd871746, 32'sd643891,
32'sd932850, 32'sd529047, 32'sd855526, 32'sd744254, 32'sd693131, 32'sd806762, 32'sd1059714, 32'sd1173052, 32'sd1180535, 32'sd976221, 32'sd845784, 32'sd516872, 32'sd1186024, 32'sd1156009,
32'sd834699, 32'sd619123, 32'sd1109172, 32'sd967433, 32'sd1151948, 32'sd922104, 32'sd578389, 32'sd404358, 32'sd652421, 32'sd586629, 32'sd660255, 32'sd858480, 32'sd1013630, 32'sd753343,
32'sd1001770, 32'sd595837, 32'sd961599, 32'sd475822, 32'sd824956, 32'sd683122, 32'sd1029490, 32'sd802134, 32'sd1114181, 32'sd604177, 32'sd992280, 32'sd1056393, 32'sd799865, 32'sd1155407,
32'sd928742, 32'sd784815, 32'sd536769, 32'sd425680, 32'sd622128, 32'sd793664, 32'sd626641, 32'sd882366, 32'sd864907, 32'sd459875, 32'sd1140007, 32'sd531854, 32'sd1051199, 32'sd532143,
32'sd1080751, 32'sd1175258, 32'sd621801, 32'sd405558, 32'sd834397, 32'sd444929, 32'sd880964, 32'sd1057345, 32'sd623216, 32'sd854115, 32'sd416953, 32'sd941217, 32'sd741353, 32'sd718964,
32'sd1107598, 32'sd787341, 32'sd773138, 32'sd1140236, 32'sd767546, 32'sd738536, 32'sd976514, 32'sd507227, 32'sd470388, 32'sd862464, 32'sd619636, 32'sd1082829, 32'sd874807, 32'sd462363,
32'sd1173554, 32'sd936340, 32'sd1021900, 32'sd589649, 32'sd854252, 32'sd1185993, 32'sd459064, 32'sd916399, 32'sd535608, 32'sd1203368, 32'sd826128, 32'sd813215, 32'sd710565, 32'sd1198160,
32'sd1167739, 32'sd891740, 32'sd537708, 32'sd553725, 32'sd771521, 32'sd891854, 32'sd710558, 32'sd527097, 32'sd911566, 32'sd431957, 32'sd595413, 32'sd893772, 32'sd543413, 32'sd643885,
32'sd562021, 32'sd618534, 32'sd940175, 32'sd1010732, 32'sd927771, 32'sd527020, 32'sd1066416, 32'sd486584, 32'sd612073, 32'sd685767, 32'sd922759, 32'sd1117590, 32'sd944725, 32'sd985961,
32'sd638939, 32'sd1178361, 32'sd461783, 32'sd796543, 32'sd482515, 32'sd770100, 32'sd1180879, 32'sd590891, 32'sd1163559, 32'sd594272, 32'sd747704, 32'sd762147, 32'sd467703, 32'sd989199,
32'sd576503, 32'sd1179643, 32'sd440171, 32'sd737166, 32'sd843471, 32'sd917850, 32'sd942637, 32'sd838563, 32'sd467290, 32'sd850328, 32'sd762514, 32'sd960770, 32'sd583897, 32'sd511047,
32'sd810537, 32'sd1065171, 32'sd684857, 32'sd414234, 32'sd635817, 32'sd409646, 32'sd1015919, 32'sd718402, 32'sd686201, 32'sd438941, 32'sd851296, 32'sd587191, 32'sd919000, 32'sd687269,
32'sd676975, 32'sd855439, 32'sd1023555, 32'sd750369, 32'sd538032, 32'sd760805, 32'sd465609, 32'sd666419, 32'sd749059, 32'sd717764, 32'sd626610, 32'sd915803, 32'sd778623, 32'sd580909,
32'sd953858, 32'sd448643, 32'sd1156296, 32'sd1077817, 32'sd666127, 32'sd497453, 32'sd499715, 32'sd443618, 32'sd589805, 32'sd511204, 32'sd1057403, 32'sd614342, 32'sd614161, 32'sd713730,
32'sd707280, 32'sd752403, 32'sd1018383, 32'sd418716, 32'sd1131629, 32'sd687853, 32'sd1172641, 32'sd664833, 32'sd1026654, 32'sd495235, 32'sd527324, 32'sd921466, 32'sd902938, 32'sd542181,
32'sd465474, 32'sd1071281, 32'sd692212, 32'sd901689, 32'sd417835, 32'sd502764, 32'sd634010, 32'sd602940, 32'sd909652, 32'sd525775, 32'sd1047641, 32'sd695407, 32'sd749410, 32'sd493992,
32'sd1197391, 32'sd447846, 32'sd518296, 32'sd659567, 32'sd741089, 32'sd987678, 32'sd930757, 32'sd839018, 32'sd565390, 32'sd857782, 32'sd1072864, 32'sd766682, 32'sd723354, 32'sd601399,
32'sd833761, 32'sd780074, 32'sd781507, 32'sd999200, 32'sd776943, 32'sd738820, 32'sd622758, 32'sd842931, 32'sd1087915, 32'sd966310, 32'sd565601, 32'sd1148868, 32'sd485584, 32'sd649436,
32'sd490573, 32'sd805088, 32'sd850138, 32'sd487062, 32'sd660434, 32'sd497581, 32'sd809115, 32'sd1201345, 32'sd947129, 32'sd1114056, 32'sd1163629, 32'sd861671, 32'sd1018203, 32'sd607426,
32'sd879085, 32'sd737895, 32'sd1177567, 32'sd955655, 32'sd921944, 32'sd639503, 32'sd1098710, 32'sd757405, 32'sd783750, 32'sd514615, 32'sd1035248, 32'sd889359, 32'sd996198, 32'sd613243,
32'sd1119957, 32'sd483679, 32'sd1200499, 32'sd1146900, 32'sd777499, 32'sd912296, 32'sd506004, 32'sd512134, 32'sd450039, 32'sd710337, 32'sd1088688, 32'sd651973, 32'sd472670, 32'sd937245,
32'sd668886, 32'sd926679, 32'sd904997, 32'sd1107550, 32'sd664959, 32'sd703524, 32'sd926357, 32'sd1010040, 32'sd1039326, 32'sd963292, 32'sd648066, 32'sd407675, 32'sd785268, 32'sd1169271,
32'sd1046124, 32'sd622817, 32'sd1100339, 32'sd787065, 32'sd513330, 32'sd606921, 32'sd1164619, 32'sd866946, 32'sd983978, 32'sd847176, 32'sd1170731, 32'sd817639, 32'sd622666, 32'sd1175498,
32'sd755302, 32'sd766632, 32'sd802984, 32'sd867734, 32'sd1046591, 32'sd485256, 32'sd1144608, 32'sd800978, 32'sd943560, 32'sd665122, 32'sd429377, 32'sd490859, 32'sd840237, 32'sd914453,
32'sd434413, 32'sd897404, 32'sd1063135, 32'sd755941, 32'sd1118325, 32'sd931985, 32'sd574358, 32'sd927990, 32'sd436147, 32'sd893984, 32'sd1035238, 32'sd649301, 32'sd938304, 32'sd1085491,
32'sd914501, 32'sd528007, 32'sd452398, 32'sd462874, 32'sd525430, 32'sd528908, 32'sd985809, 32'sd742800, 32'sd614442, 32'sd414026, 32'sd1164501, 32'sd1018982, 32'sd1060333, 32'sd506841,
32'sd844783, 32'sd937673, 32'sd678479, 32'sd884606, 32'sd1097923, 32'sd1053608, 32'sd1014369, 32'sd851960, 32'sd1130405, 32'sd1198660, 32'sd1048174, 32'sd616569, 32'sd1012928, 32'sd524421,
32'sd1044860, 32'sd723399, 32'sd760655, 32'sd532797, 32'sd957716, 32'sd1037148, 32'sd433753, 32'sd875710, 32'sd949656, 32'sd839924, 32'sd789383, 32'sd1148561, 32'sd835427, 32'sd793413,
32'sd504313, 32'sd767739, 32'sd496472, 32'sd982091, 32'sd1192137, 32'sd981960, 32'sd901504, 32'sd1030739, 32'sd696173, 32'sd841957, 32'sd535615, 32'sd439132, 32'sd474295, 32'sd1176346,
32'sd1024322, 32'sd1051950, 32'sd931897, 32'sd423734, 32'sd461869, 32'sd564927, 32'sd1003077, 32'sd779327, 32'sd773662, 32'sd982306, 32'sd416906, 32'sd971306, 32'sd798783, 32'sd700918,
32'sd1017602, 32'sd952083, 32'sd1176838, 32'sd1202924, 32'sd659779, 32'sd1171285, 32'sd444645, 32'sd687579, 32'sd527144, 32'sd1017658, 32'sd1134372, 32'sd1128886, 32'sd542392, 32'sd629442,
32'sd781764, 32'sd791668, 32'sd441350, 32'sd1107323, 32'sd844592, 32'sd1106419, 32'sd620004, 32'sd468926, 32'sd648807, 32'sd1028208, 32'sd906143, 32'sd773655, 32'sd870218, 32'sd811120,
32'sd715560, 32'sd786906, 32'sd995618, 32'sd794410, 32'sd809448, 32'sd498728, 32'sd636210, 32'sd773483, 32'sd975876, 32'sd593817, 32'sd1018852, 32'sd943322, 32'sd1139047, 32'sd587931,
32'sd597930, 32'sd454016, 32'sd1102066, 32'sd992160, 32'sd515358, 32'sd1066573, 32'sd608759, 32'sd563450, 32'sd768538, 32'sd1203277, 32'sd513477, 32'sd438617, 32'sd800827, 32'sd698729,
32'sd684268, 32'sd859168, 32'sd515642, 32'sd556783, 32'sd624451, 32'sd686760, 32'sd855947, 32'sd1045587, 32'sd1143875, 32'sd910089, 32'sd487008, 32'sd916916, 32'sd892020, 32'sd483911,
32'sd1002816, 32'sd606276, 32'sd566424, 32'sd817435, 32'sd1115649, 32'sd625976, 32'sd753856, 32'sd1193033, 32'sd679796, 32'sd575378, 32'sd915346, 32'sd608254, 32'sd787125, 32'sd1138340,
32'sd616169, 32'sd418343, 32'sd612660, 32'sd975764, 32'sd426875, 32'sd1150164, 32'sd961747, 32'sd919852, 32'sd1013010, 32'sd756520, 32'sd816795, 32'sd1142467, 32'sd571519, 32'sd651476,
32'sd1057464, 32'sd407124, 32'sd549707, 32'sd516701, 32'sd667969, 32'sd678730, 32'sd1115893, 32'sd875296, 32'sd749972, 32'sd729475, 32'sd789823, 32'sd1058339, 32'sd568599, 32'sd1160757,
32'sd1001011, 32'sd423817, 32'sd660838, 32'sd1119204, 32'sd505015, 32'sd552174, 32'sd1205108, 32'sd900938, 32'sd790892, 32'sd435571, 32'sd996119, 32'sd1047685, 32'sd485259, 32'sd736747,
32'sd1135409, 32'sd682048, 32'sd516104, 32'sd492568, 32'sd757515, 32'sd815623, 32'sd867720, 32'sd703607, 32'sd444967, 32'sd482560, 32'sd890961, 32'sd819250, 32'sd1181122, 32'sd819306,
32'sd958308, 32'sd539838, 32'sd1163320, 32'sd443958, 32'sd630636, 32'sd1202150, 32'sd556585, 32'sd1108091, 32'sd541436, 32'sd720403, 32'sd623676, 32'sd540785, 32'sd537790, 32'sd900014,
32'sd569506, 32'sd446969, 32'sd863223, 32'sd569020, 32'sd1116456, 32'sd1095819, 32'sd506290, 32'sd1044302, 32'sd442442, 32'sd520410, 32'sd885516, 32'sd1069186, 32'sd483060, 32'sd1078087,
32'sd898345, 32'sd902542, 32'sd898920, 32'sd523135, 32'sd903817, 32'sd796743, 32'sd1154088, 32'sd1128755, 32'sd642679, 32'sd1062907, 32'sd843456, 32'sd803562, 32'sd865154, 32'sd795411,
32'sd1209222, 32'sd727481, 32'sd517395, 32'sd832387, 32'sd1045209, 32'sd455973, 32'sd1208961, 32'sd1062060, 32'sd470310, 32'sd860528, 32'sd684295, 32'sd465696, 32'sd717346, 32'sd460039,
32'sd651820, 32'sd1148764, 32'sd775011, 32'sd776930, 32'sd887612, 32'sd442914, 32'sd1120956, 32'sd625861, 32'sd788637, 32'sd747616, 32'sd462950, 32'sd707810, 32'sd1011722, 32'sd1021137,
32'sd571967, 32'sd1139647, 32'sd641530, 32'sd939149, 32'sd751974, 32'sd618190, 32'sd480242, 32'sd470682, 32'sd1059521, 32'sd612836, 32'sd823587, 32'sd543914, 32'sd730594, 32'sd789178,
32'sd624728, 32'sd476413, 32'sd455266, 32'sd1196634, 32'sd858688, 32'sd763094, 32'sd810497, 32'sd877639, 32'sd569213, 32'sd639704, 32'sd1197799, 32'sd736090, 32'sd743831, 32'sd535896,
32'sd996042, 32'sd575568, 32'sd1054771, 32'sd794997, 32'sd723376, 32'sd864114, 32'sd880456, 32'sd783109, 32'sd683851, 32'sd1029968, 32'sd988090, 32'sd867091, 32'sd898153, 32'sd1004434,
32'sd1003773, 32'sd651924, 32'sd963852, 32'sd882915, 32'sd1056375, 32'sd1127565, 32'sd467695, 32'sd511731, 32'sd690425, 32'sd589604, 32'sd729284, 32'sd1026036, 32'sd1025108, 32'sd896634,
32'sd487586, 32'sd541691, 32'sd506364, 32'sd480232, 32'sd1095756, 32'sd1112684, 32'sd941742, 32'sd674169, 32'sd878081, 32'sd1032458, 32'sd490308, 32'sd895566, 32'sd1174693, 32'sd713913,
32'sd1159905, 32'sd591643, 32'sd623565, 32'sd440529, 32'sd1111853, 32'sd847924, 32'sd727932, 32'sd895941, 32'sd973557, 32'sd884811, 32'sd611088, 32'sd604163, 32'sd887508, 32'sd425033,
32'sd553882, 32'sd1035871, 32'sd1025114, 32'sd666641, 32'sd416687, 32'sd1034314, 32'sd481842, 32'sd703758, 32'sd726769, 32'sd1111571, 32'sd565456, 32'sd1107346, 32'sd590557, 32'sd1178023,
32'sd661541, 32'sd1055596, 32'sd905134, 32'sd1132387, 32'sd535108, 32'sd1168532, 32'sd693101, 32'sd668274, 32'sd774921, 32'sd1072038, 32'sd1170082, 32'sd968719, 32'sd718453, 32'sd1007748,
32'sd432871, 32'sd510050, 32'sd875248, 32'sd548482, 32'sd702368, 32'sd1083301, 32'sd724489, 32'sd712082, 32'sd564366, 32'sd584460, 32'sd843296, 32'sd595910, 32'sd924527, 32'sd868950,
32'sd957167, 32'sd499036, 32'sd616046, 32'sd872378, 32'sd406069, 32'sd829459, 32'sd587553, 32'sd933146, 32'sd788544, 32'sd867029, 32'sd1079264, 32'sd431199, 32'sd482563, 32'sd529551,
32'sd905250, 32'sd861366, 32'sd596762, 32'sd1141542, 32'sd835092, 32'sd933794, 32'sd688017, 32'sd737822, 32'sd988168, 32'sd445092, 32'sd581099, 32'sd734648, 32'sd528332, 32'sd1040594,
32'sd1020399, 32'sd1134832, 32'sd1035592, 32'sd928743, 32'sd970241, 32'sd808937, 32'sd466572, 32'sd1103197, 32'sd537433, 32'sd582186, 32'sd784220, 32'sd709896, 32'sd1015317, 32'sd653127,
32'sd621586, 32'sd909461, 32'sd611412, 32'sd1183190, 32'sd657480, 32'sd943648, 32'sd862505, 32'sd472091, 32'sd913913, 32'sd594627, 32'sd1052597, 32'sd1096550, 32'sd906304, 32'sd868362,
32'sd640098, 32'sd660141, 32'sd550745, 32'sd678667, 32'sd702259, 32'sd993377, 32'sd591801, 32'sd795641, 32'sd1121654, 32'sd617524, 32'sd1116368, 32'sd1082579, 32'sd924122, 32'sd485770,
32'sd957997, 32'sd445635, 32'sd672370, 32'sd773245, 32'sd458880, 32'sd1032409, 32'sd1083379, 32'sd1040660, 32'sd863981, 32'sd933442, 32'sd1004114, 32'sd840500, 32'sd686396, 32'sd843919,
32'sd794538, 32'sd503893, 32'sd919201, 32'sd612129, 32'sd1164553, 32'sd1004810, 32'sd595562, 32'sd1074498, 32'sd805100, 32'sd861603, 32'sd591591, 32'sd767002, 32'sd699579, 32'sd826925,
32'sd1128382, 32'sd947413, 32'sd849596, 32'sd808553, 32'sd542477, 32'sd1106731, 32'sd1188566, 32'sd893741, 32'sd870219, 32'sd726262, 32'sd811502, 32'sd776520, 32'sd1013046, 32'sd1185370,
32'sd946035, 32'sd410435, 32'sd411889, 32'sd815884, 32'sd1050294, 32'sd407384, 32'sd597499, 32'sd720482, 32'sd605609, 32'sd929992, 32'sd679045, 32'sd710774, 32'sd805593, 32'sd554538,
32'sd736505, 32'sd699992, 32'sd469509, 32'sd683123, 32'sd453814, 32'sd1118246, 32'sd462468, 32'sd674646, 32'sd523068, 32'sd599190, 32'sd967859, 32'sd509606, 32'sd1122232, 32'sd960451,
32'sd523391, 32'sd572310, 32'sd851601, 32'sd667055, 32'sd1186341, 32'sd749168, 32'sd838829, 32'sd659517, 32'sd1000130, 32'sd618188, 32'sd415297, 32'sd754180, 32'sd879810, 32'sd726554,
32'sd707934, 32'sd1168060, 32'sd854217, 32'sd705044, 32'sd932891, 32'sd753301, 32'sd529523, 32'sd941283, 32'sd530410, 32'sd1206598, 32'sd1137333, 32'sd558427, 32'sd867538, 32'sd1024489,
32'sd1043901, 32'sd499022, 32'sd1073779, 32'sd721878, 32'sd843374, 32'sd757632, 32'sd623088, 32'sd528601, 32'sd1074026, 32'sd523078, 32'sd831698, 32'sd834679, 32'sd1107933, 32'sd981556,
32'sd724599, 32'sd799606, 32'sd1036052, 32'sd1113689, 32'sd485587, 32'sd1056803, 32'sd875270, 32'sd1050839, 32'sd861053, 32'sd698819, 32'sd584736, 32'sd745413, 32'sd513838, 32'sd1102233,
32'sd806415, 32'sd1113354, 32'sd1125782, 32'sd734731, 32'sd867139, 32'sd484746, 32'sd513526, 32'sd1025987, 32'sd813937, 32'sd800601, 32'sd1152752, 32'sd409997, 32'sd637640, 32'sd623338,
32'sd1173596, 32'sd404944, 32'sd518917, 32'sd535639, 32'sd627636, 32'sd945280, 32'sd490301, 32'sd832350, 32'sd984408, 32'sd613232, 32'sd796868, 32'sd688781, 32'sd1111445, 32'sd1176425,
32'sd640699, 32'sd959003, 32'sd1100888, 32'sd446524, 32'sd410313, 32'sd1062275, 32'sd767717, 32'sd990013, 32'sd1191888, 32'sd448223, 32'sd1130599, 32'sd475512, 32'sd627003, 32'sd1102407,
32'sd785732, 32'sd1182604, 32'sd702590, 32'sd1049728, 32'sd419280, 32'sd561943, 32'sd610392, 32'sd831220, 32'sd593800, 32'sd1184315, 32'sd780557, 32'sd573343, 32'sd1143897, 32'sd587621,
32'sd923380, 32'sd456805, 32'sd733470, 32'sd523163, 32'sd694787, 32'sd994582, 32'sd412440, 32'sd843005, 32'sd864692, 32'sd489319, 32'sd466542, 32'sd768958, 32'sd723712, 32'sd1195132,
32'sd886495, 32'sd588053, 32'sd863028, 32'sd1197704, 32'sd819665, 32'sd523701, 32'sd537867, 32'sd494376, 32'sd1111236, 32'sd519810, 32'sd559209, 32'sd922529, 32'sd560487, 32'sd1046664,
32'sd895447, 32'sd705793, 32'sd657522, 32'sd492824, 32'sd627186, 32'sd1148859, 32'sd536805, 32'sd558229, 32'sd1208346, 32'sd1149817, 32'sd1060774, 32'sd750734, 32'sd517948, 32'sd892460,
32'sd601979, 32'sd1157159, 32'sd448742, 32'sd800775, 32'sd836561, 32'sd1103063, 32'sd1152743, 32'sd439435, 32'sd555265, 32'sd425755, 32'sd740915, 32'sd842348, 32'sd871062, 32'sd714850,
32'sd816989, 32'sd1004051, 32'sd956338, 32'sd469984, 32'sd783809, 32'sd1058402, 32'sd562068, 32'sd857503, 32'sd786783, 32'sd506171, 32'sd1022825, 32'sd605812, 32'sd1062337, 32'sd1166138,
32'sd684078, 32'sd808672, 32'sd690140, 32'sd737492, 32'sd447351, 32'sd1154374, 32'sd562575, 32'sd850726, 32'sd1164301, 32'sd573842, 32'sd846946, 32'sd1093752, 32'sd1175651, 32'sd890040

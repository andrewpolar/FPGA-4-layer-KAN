32'sd133861, 32'sd77671, 32'sd50580, 32'sd245928, 32'sd296976, 32'sd1031824, 32'sd240636, 32'sd361405, 32'sd522667, 32'sd520401,
32'sd9048, 32'sd58582, 32'sd155186, 32'sd87153, 32'sd681627, 32'sd756133, 32'sd563715, 32'sd518132, 32'sd192813, 32'sd242749,
32'sd266116, 32'sd106352, 32'sd29422, 32'sd34802, 32'sd224613, 32'sd207739, 32'sd242616, 32'sd396466, 32'sd207819, 32'sd57132,
32'sd381798, 32'sd627443, 32'sd244538, 32'sd50979, 32'sd272052, 32'sd81971, 32'sd196878, 32'sd61654, 32'sd61959, 32'sd333791,
32'sd51432, 32'sd1086353, 32'sd311934, 32'sd189225, 32'sd14148, 32'sd438228, 32'sd7741, 32'sd304247, 32'sd269955, 32'sd408246,
32'sd826567, 32'sd86836, 32'sd173742, 32'sd16234, 32'sd516954, 32'sd280130, 32'sd292696, 32'sd82927, 32'sd154398, 32'sd977292,
32'sd142654, 32'sd667025, 32'sd471152, 32'sd68433, 32'sd153216, 32'sd176450, 32'sd271124, 32'sd24024, 32'sd322356, 32'sd466471,
32'sd636505, 32'sd403815, 32'sd448934, 32'sd223196, 32'sd34792, 32'sd20452, 32'sd174484, 32'sd277057, 32'sd365954, 32'sd292492,
32'sd24661, 32'sd38909, 32'sd314686, 32'sd1016058, 32'sd372933, 32'sd373551, 32'sd257418, 32'sd10470, 32'sd431964, 32'sd63742,
32'sd161604, 32'sd142772, 32'sd61770, 32'sd367993, 32'sd17944, 32'sd4281, 32'sd72244, 32'sd144570, 32'sd160599, 32'sd6485,
32'sd170714, 32'sd123246, 32'sd245491, 32'sd189984, 32'sd67097, 32'sd92823, 32'sd84877, 32'sd444558, 32'sd315455, 32'sd161307,
32'sd498067, 32'sd272185, 32'sd270186, 32'sd45173, 32'sd269333, 32'sd81106, 32'sd106578, 32'sd1244002, 32'sd409648, 32'sd42316,
32'sd40466, 32'sd527692, 32'sd284836, 32'sd886099, 32'sd266903, 32'sd130428, 32'sd521619, 32'sd690430, 32'sd244453, 32'sd28018,
32'sd142283, 32'sd351207, 32'sd598134, 32'sd284117, 32'sd520394, 32'sd151992, 32'sd406976, 32'sd139615, 32'sd330062, 32'sd177735,
32'sd347105, 32'sd117852, 32'sd103366, 32'sd204004, 32'sd204422, 32'sd149679, 32'sd6437, 32'sd104706, 32'sd267066, 32'sd603268,
32'sd778708, 32'sd13482, 32'sd177798, 32'sd545806, 32'sd471299, 32'sd552594, 32'sd180775, 32'sd505003, 32'sd666690, 32'sd31906,
32'sd96102, 32'sd1058663, 32'sd382380, 32'sd443802, 32'sd21939, 32'sd747036, 32'sd316690, 32'sd184895, 32'sd127984, 32'sd132413,
32'sd100816, 32'sd690657, 32'sd219594, 32'sd846251, 32'sd182684, 32'sd31635, 32'sd214740, 32'sd68236, 32'sd2296, 32'sd21699,
32'sd138699, 32'sd134382, 32'sd107205, 32'sd262, 32'sd5408, 32'sd151236, 32'sd112124, 32'sd146230, 32'sd87923, 32'sd321069,
32'sd70359, 32'sd84410, 32'sd383680, 32'sd325135, 32'sd58452, 32'sd19578, 32'sd519890, 32'sd462006, 32'sd617640, 32'sd21029,
32'sd121542, 32'sd187129, 32'sd84222, 32'sd152758, 32'sd265862, 32'sd201514, 32'sd6901, 32'sd235667, 32'sd240704, 32'sd122877,
32'sd164915, 32'sd360483, 32'sd190499, 32'sd202062, 32'sd52453, 32'sd217508, 32'sd212593, 32'sd83215, 32'sd528948, 32'sd26631,
32'sd90730, 32'sd730923, 32'sd265343, 32'sd156016, 32'sd188482, 32'sd574410, 32'sd93829, 32'sd623919, 32'sd264157, 32'sd418170,
32'sd536916, 32'sd365500, 32'sd186489, 32'sd331128, 32'sd494966, 32'sd283816, 32'sd133556, 32'sd284439, 32'sd122692, 32'sd250601,
32'sd231649, 32'sd468591, 32'sd53352, 32'sd311069, 32'sd420791, 32'sd1281159, 32'sd117124, 32'sd89677, 32'sd82204, 32'sd52613,
32'sd18980, 32'sd306932, 32'sd386032, 32'sd24129, 32'sd276734, 32'sd263377, 32'sd280566, 32'sd334863, 32'sd194267, 32'sd717781,
32'sd344562, 32'sd197670, 32'sd140195, 32'sd1049531, 32'sd287782, 32'sd35348, 32'sd827253, 32'sd161274, 32'sd186958, 32'sd432839,
32'sd298694, 32'sd200636, 32'sd591899, 32'sd473370, 32'sd416623, 32'sd471871, 32'sd109808, 32'sd140116, 32'sd553905, 32'sd495957,
32'sd380265, 32'sd463353, 32'sd18119, 32'sd304025, 32'sd233697, 32'sd440765, 32'sd138605, 32'sd836915, 32'sd420970, 32'sd271009,
32'sd508890, 32'sd202600, 32'sd471792, 32'sd43931, 32'sd162806, 32'sd47291, 32'sd100599, 32'sd53227, 32'sd105338, 32'sd368111,
32'sd555513, 32'sd79160, 32'sd61649, 32'sd54031, 32'sd73309, 32'sd628526, 32'sd687053, 32'sd3933, 32'sd215220, 32'sd871498,
32'sd872805, 32'sd619097, 32'sd423088, 32'sd2876, 32'sd349105, 32'sd221406, 32'sd247572, 32'sd4137, 32'sd292042, 32'sd77988,
32'sd86375, 32'sd144072, 32'sd243073, 32'sd4345, 32'sd29406, 32'sd23468, 32'sd87072, 32'sd309401, 32'sd183185, 32'sd265402,
32'sd168011, 32'sd102263, 32'sd550074, 32'sd237458, 32'sd16538, 32'sd14580, 32'sd257324, 32'sd264954, 32'sd213023, 32'sd39559,
32'sd136166, 32'sd378779, 32'sd6139, 32'sd87279, 32'sd78273, 32'sd181300, 32'sd63069, 32'sd698241, 32'sd272952, 32'sd566506,
32'sd529179, 32'sd104991, 32'sd211242, 32'sd83296, 32'sd128402, 32'sd709176, 32'sd216812, 32'sd18373, 32'sd480170, 32'sd157708,
32'sd622331, 32'sd367431, 32'sd128715, 32'sd231390, 32'sd631244, 32'sd726051, 32'sd5023, 32'sd1424, 32'sd344570, 32'sd146634,
32'sd300185, 32'sd331104, 32'sd591723, 32'sd267330, 32'sd492438, 32'sd291825, 32'sd330209, 32'sd116695, 32'sd35736, 32'sd13237,
32'sd620841, 32'sd603000, 32'sd73742, 32'sd509953, 32'sd10320, 32'sd413905, 32'sd451765, 32'sd115147, 32'sd205543, 32'sd55069,
32'sd505871, 32'sd29073, 32'sd230669, 32'sd421434, 32'sd817209, 32'sd314048, 32'sd777359, 32'sd87549, 32'sd962199, 32'sd381633,
32'sd348381, 32'sd57922, 32'sd258065, 32'sd178342, 32'sd91847, 32'sd88104, 32'sd445191, 32'sd46510, 32'sd191601, 32'sd182604,
32'sd94223, 32'sd30562, 32'sd281103, 32'sd600844, 32'sd127406, 32'sd209837, 32'sd389272, 32'sd1223377, 32'sd328558, 32'sd18294,
32'sd315392, 32'sd150943, 32'sd788648, 32'sd251364, 32'sd437656, 32'sd478927, 32'sd685596, 32'sd100713, 32'sd303860, 32'sd213089,
32'sd614761, 32'sd208297, 32'sd318648, 32'sd691479, 32'sd106457, 32'sd6697, 32'sd1430, 32'sd144221, 32'sd145128, 32'sd54279,
32'sd145659, 32'sd561429, 32'sd222146, 32'sd107533, 32'sd381518, 32'sd211496, 32'sd470984, 32'sd309660, 32'sd135285, 32'sd175027,
32'sd418577, 32'sd9606, 32'sd564030, 32'sd90800, 32'sd350071, 32'sd335522, 32'sd141841, 32'sd618364, 32'sd760744, 32'sd278769,
32'sd395597, 32'sd52524, 32'sd256557, 32'sd217402, 32'sd298950, 32'sd327296, 32'sd181783, 32'sd31672, 32'sd396410, 32'sd942954,
32'sd133213, 32'sd124649, 32'sd169016, 32'sd202644, 32'sd46970, 32'sd28564, 32'sd398175, 32'sd47170, 32'sd234293, 32'sd241849,
32'sd200731, 32'sd872293, 32'sd334095, 32'sd108299, 32'sd1169268, 32'sd275670, 32'sd198978, 32'sd251869, 32'sd476022, 32'sd76442,
32'sd35241, 32'sd84145, 32'sd443785, 32'sd570424, 32'sd66323, 32'sd336679, 32'sd54840, 32'sd102632, 32'sd803270, 32'sd26099,
32'sd294845, 32'sd214113, 32'sd663710, 32'sd297999, 32'sd31063, 32'sd556976, 32'sd30801, 32'sd173541, 32'sd133731, 32'sd393094,
32'sd364469, 32'sd420609, 32'sd200090, 32'sd126299, 32'sd189607, 32'sd110433, 32'sd351357, 32'sd99973, 32'sd166536, 32'sd507885,
32'sd158325, 32'sd106290, 32'sd389007, 32'sd3601, 32'sd87084, 32'sd1017937, 32'sd575314, 32'sd417456, 32'sd140944, 32'sd336931,
32'sd206279, 32'sd48252, 32'sd220426, 32'sd188363, 32'sd230463, 32'sd232639, 32'sd959483, 32'sd331006, 32'sd199119, 32'sd60875,
32'sd83406, 32'sd238580, 32'sd186395, 32'sd21540, 32'sd29091, 32'sd234142, 32'sd442613, 32'sd360975, 32'sd107822, 32'sd904654,
32'sd650547, 32'sd233816, 32'sd35149, 32'sd102874, 32'sd210624, 32'sd722978, 32'sd523412, 32'sd220570, 32'sd113838, 32'sd278277,
32'sd307801, 32'sd262520, 32'sd194486, 32'sd131158, 32'sd196189, 32'sd169785, 32'sd329352, 32'sd183583, 32'sd41107, 32'sd453568,
32'sd57987, 32'sd204918, 32'sd258882, 32'sd68154, 32'sd148894, 32'sd163996, 32'sd821254, 32'sd307, 32'sd361126, 32'sd60029,
32'sd4625, 32'sd239664, 32'sd442083, 32'sd267921, 32'sd40357, 32'sd361768, 32'sd1130698, 32'sd324081, 32'sd137207, 32'sd373596,
32'sd478695, 32'sd144749, 32'sd93585, 32'sd912234, 32'sd691061, 32'sd51583, 32'sd103926, 32'sd32811, 32'sd263010, 32'sd323977,
32'sd257584, 32'sd404792, 32'sd61505, 32'sd501077, 32'sd277626, 32'sd481312, 32'sd128794, 32'sd663464, 32'sd464506, 32'sd283895,
32'sd33565, 32'sd161459, 32'sd99982, 32'sd541861, 32'sd243975, 32'sd135038, 32'sd429949, 32'sd332263, 32'sd261945, 32'sd747765,
32'sd270217, 32'sd727077, 32'sd119377, 32'sd859122, 32'sd403531, 32'sd129060, 32'sd71716, 32'sd481192, 32'sd89320, 32'sd645138,
32'sd337418, 32'sd121562, 32'sd145430, 32'sd367825, 32'sd543124, 32'sd193337, 32'sd65344, 32'sd567833, 32'sd370533, 32'sd234132,
32'sd271311, 32'sd2836, 32'sd58675, 32'sd438717, 32'sd29680, 32'sd4569, 32'sd359298, 32'sd1224964, 32'sd782414, 32'sd34788,
32'sd204820, 32'sd89120, 32'sd481610, 32'sd395703, 32'sd96162, 32'sd418124, 32'sd391740, 32'sd292932, 32'sd1027542, 32'sd46942,
32'sd81795, 32'sd150900, 32'sd964411, 32'sd61679, 32'sd810591, 32'sd30859, 32'sd418157, 32'sd26867, 32'sd47202, 32'sd174816,
32'sd183298, 32'sd240774, 32'sd433022, 32'sd380255, 32'sd753043, 32'sd64572, 32'sd294, 32'sd196273, 32'sd80257, 32'sd56884,
32'sd259037, 32'sd35899, 32'sd168561, 32'sd551726, 32'sd589392, 32'sd563186, 32'sd441660, 32'sd408304, 32'sd10492, 32'sd55516,
32'sd192367, 32'sd403088, 32'sd568011, 32'sd47617, 32'sd18963, 32'sd602384, 32'sd440272, 32'sd45546, 32'sd143464, 32'sd209512,
32'sd93182, 32'sd159246, 32'sd384340, 32'sd611308, 32'sd10024, 32'sd873135, 32'sd219950, 32'sd63108, 32'sd387816, 32'sd775825,
32'sd254665, 32'sd568026, 32'sd7325, 32'sd611581, 32'sd85300, 32'sd137802, 32'sd245716, 32'sd431394, 32'sd116101, 32'sd1094568,
32'sd8878, 32'sd1025876, 32'sd1063120, 32'sd440123, 32'sd117189, 32'sd241366, 32'sd93503, 32'sd141517, 32'sd235750, 32'sd118943,
32'sd15897, 32'sd708107, 32'sd236905, 32'sd149735, 32'sd518372, 32'sd898644, 32'sd65484, 32'sd224049, 32'sd332608, 32'sd176109,
32'sd168742, 32'sd177196, 32'sd180684, 32'sd209776, 32'sd402387, 32'sd29029, 32'sd30916, 32'sd228772, 32'sd38920, 32'sd146667,
32'sd426484, 32'sd327740, 32'sd101420, 32'sd1180797, 32'sd460031, 32'sd140170, 32'sd256999, 32'sd63688, 32'sd653031, 32'sd502149,
32'sd70092, 32'sd440591, 32'sd359940, 32'sd207852, 32'sd418395, 32'sd235222, 32'sd761808, 32'sd220829, 32'sd103972, 32'sd181717,
32'sd461456, 32'sd58086, 32'sd1110389, 32'sd103768, 32'sd342283, 32'sd171209, 32'sd13058, 32'sd486162, 32'sd572897, 32'sd398249,
32'sd197744, 32'sd6035, 32'sd554500, 32'sd30293, 32'sd536084, 32'sd1004074, 32'sd725145, 32'sd576955, 32'sd379775, 32'sd569428,
32'sd290837, 32'sd209495, 32'sd80040, 32'sd55506, 32'sd376757, 32'sd19321, 32'sd168667, 32'sd13917, 32'sd8446, 32'sd496294,
32'sd29775, 32'sd24701, 32'sd610892, 32'sd24658, 32'sd126500, 32'sd473295, 32'sd543504, 32'sd461648, 32'sd341551, 32'sd92119,
32'sd581506, 32'sd157983, 32'sd248990, 32'sd17303, 32'sd126905, 32'sd464946, 32'sd634246, 32'sd147597, 32'sd633152, 32'sd263827,
32'sd557284, 32'sd496593, 32'sd129108, 32'sd149950, 32'sd223402, 32'sd468150, 32'sd222374, 32'sd441418, 32'sd421246, 32'sd324810,
32'sd640926, 32'sd113742, 32'sd768111, 32'sd325306, 32'sd770384, 32'sd219898, 32'sd70296, 32'sd63511, 32'sd143325, 32'sd189401,
32'sd482907, 32'sd483783, 32'sd334257, 32'sd112811, 32'sd294346, 32'sd13456, 32'sd196686, 32'sd496060, 32'sd90620, 32'sd12424,
32'sd255253, 32'sd420042, 32'sd387555, 32'sd306439, 32'sd943145, 32'sd417056, 32'sd594409, 32'sd120894, 32'sd215707, 32'sd518947,
32'sd22097, 32'sd111771, 32'sd744310, 32'sd423441, 32'sd184425, 32'sd3346, 32'sd554385, 32'sd479359, 32'sd77177, 32'sd601834,
32'sd1056480, 32'sd129337, 32'sd740065, 32'sd542699, 32'sd121674, 32'sd25449, 32'sd262, 32'sd828985, 32'sd55842, 32'sd450374,
32'sd287244, 32'sd20443, 32'sd12090, 32'sd809485, 32'sd15749, 32'sd380371, 32'sd606437, 32'sd11865, 32'sd518920, 32'sd600201,
32'sd561510, 32'sd33892, 32'sd177656, 32'sd661224, 32'sd60161, 32'sd470834, 32'sd12247, 32'sd53057, 32'sd730574, 32'sd381782,
32'sd106392, 32'sd394473, 32'sd182936, 32'sd230068, 32'sd94214, 32'sd472252, 32'sd279350, 32'sd573042, 32'sd351903, 32'sd529428,
32'sd119850, 32'sd787456, 32'sd656013, 32'sd742464, 32'sd102764, 32'sd29575, 32'sd20554, 32'sd236838, 32'sd210255, 32'sd377848,
32'sd17145, 32'sd204506, 32'sd212175, 32'sd730572, 32'sd36394, 32'sd791277, 32'sd313322, 32'sd36115, 32'sd506084, 32'sd294606,
32'sd829948, 32'sd535414, 32'sd342049, 32'sd72889, 32'sd383514, 32'sd547198, 32'sd30892, 32'sd128402, 32'sd161658, 32'sd399628,
32'sd31484, 32'sd326657, 32'sd8143, 32'sd121540, 32'sd302008, 32'sd56551, 32'sd65493, 32'sd25592, 32'sd851182, 32'sd39001,
32'sd710885, 32'sd97266, 32'sd138176, 32'sd207640, 32'sd118470, 32'sd268059, 32'sd230700, 32'sd27252, 32'sd179309, 32'sd8294,
32'sd487122, 32'sd214249, 32'sd1005822, 32'sd271291, 32'sd806625, 32'sd96837, 32'sd177960, 32'sd285307, 32'sd388920, 32'sd163360,
32'sd30551, 32'sd4641, 32'sd374548, 32'sd296631, 32'sd131671, 32'sd80288, 32'sd21667, 32'sd95383, 32'sd148888, 32'sd216686,
32'sd246250, 32'sd331043, 32'sd492928, 32'sd55391, 32'sd73032, 32'sd137370, 32'sd311971, 32'sd88694, 32'sd35373, 32'sd61639,
32'sd11266, 32'sd494727, 32'sd98681, 32'sd78936, 32'sd113897, 32'sd67157, 32'sd414964, 32'sd12306, 32'sd476765, 32'sd368836,
32'sd121554, 32'sd349773, 32'sd100718, 32'sd321382, 32'sd160433, 32'sd566467, 32'sd232890, 32'sd158777, 32'sd278233, 32'sd579664,
32'sd324194, 32'sd308860, 32'sd46471, 32'sd284956, 32'sd545046, 32'sd345282, 32'sd238408, 32'sd402420, 32'sd56699, 32'sd38066,
32'sd238376, 32'sd60456, 32'sd155856, 32'sd160468, 32'sd558103, 32'sd168789, 32'sd127812, 32'sd92863, 32'sd149941, 32'sd181225,
32'sd612216, 32'sd216812, 32'sd82284, 32'sd456196, 32'sd81840, 32'sd371365, 32'sd194833, 32'sd80118, 32'sd66667, 32'sd186349,
32'sd136220, 32'sd174910, 32'sd314483, 32'sd522525, 32'sd29578, 32'sd547473, 32'sd129078, 32'sd326163, 32'sd19368, 32'sd17405,
32'sd209966, 32'sd219102, 32'sd175345, 32'sd343420, 32'sd264415, 32'sd144928, 32'sd633584, 32'sd228728, 32'sd213715, 32'sd43206,
32'sd1074595, 32'sd574518, 32'sd129908, 32'sd234756, 32'sd253429, 32'sd505541, 32'sd314355, 32'sd19731, 32'sd304226, 32'sd235017,
32'sd334989, 32'sd310312, 32'sd18868, 32'sd111954, 32'sd118425, 32'sd704114, 32'sd188541, 32'sd168196, 32'sd3234, 32'sd316115,
32'sd196352, 32'sd18594, 32'sd11398, 32'sd163862, 32'sd305425, 32'sd429417, 32'sd881239, 32'sd25327, 32'sd462358, 32'sd73316,
32'sd69847, 32'sd225948, 32'sd107467, 32'sd886460, 32'sd210327, 32'sd129354, 32'sd95442, 32'sd55822, 32'sd243531, 32'sd235557,
32'sd355495, 32'sd295761, 32'sd33846, 32'sd110949, 32'sd69148, 32'sd1137188, 32'sd118377, 32'sd400450, 32'sd6732, 32'sd380680,
32'sd30569, 32'sd46660, 32'sd108364, 32'sd3067, 32'sd90349, 32'sd17133, 32'sd91007, 32'sd210204, 32'sd377191, 32'sd684594,
32'sd27675, 32'sd229727, 32'sd171546, 32'sd308350, 32'sd386863, 32'sd61707, 32'sd142980, 32'sd484512, 32'sd223239, 32'sd242711,
32'sd299029, 32'sd120220, 32'sd614487, 32'sd134225, 32'sd32936, 32'sd213626, 32'sd25422, 32'sd90987, 32'sd357083, 32'sd381508,
32'sd86416, 32'sd1296204, 32'sd394380, 32'sd751975, 32'sd51838, 32'sd612103, 32'sd47519, 32'sd1001926, 32'sd194039, 32'sd22985,
32'sd158774, 32'sd544152, 32'sd1297563, 32'sd76977, 32'sd153751, 32'sd63414, 32'sd318356, 32'sd809002, 32'sd644832, 32'sd280827,
32'sd681830, 32'sd26915, 32'sd39111, 32'sd594531, 32'sd105421, 32'sd534973, 32'sd147004, 32'sd264445, 32'sd161824, 32'sd66572,
32'sd50290, 32'sd79878, 32'sd516966, 32'sd53541, 32'sd494868, 32'sd425500, 32'sd278711, 32'sd21238, 32'sd401908, 32'sd249250,
32'sd69771, 32'sd224494, 32'sd167666, 32'sd152045, 32'sd42619, 32'sd379746, 32'sd535665, 32'sd360919, 32'sd159092, 32'sd107852,
32'sd115176, 32'sd308281, 32'sd63708, 32'sd679360, 32'sd12399, 32'sd692520, 32'sd14063, 32'sd664223, 32'sd141925, 32'sd377335,
32'sd391698, 32'sd464960, 32'sd135071, 32'sd96470, 32'sd656442, 32'sd25674, 32'sd85376, 32'sd11646, 32'sd1116645, 32'sd77271,
32'sd81357, 32'sd241116, 32'sd1121284, 32'sd393250, 32'sd212655, 32'sd368425, 32'sd397352, 32'sd254127, 32'sd838938, 32'sd212764,
32'sd686080, 32'sd1100155, 32'sd535175, 32'sd749528, 32'sd84723, 32'sd127321, 32'sd713135, 32'sd13877, 32'sd173769, 32'sd31545,
32'sd788449, 32'sd210291, 32'sd459041, 32'sd762384, 32'sd97479, 32'sd154074, 32'sd303196, 32'sd351676, 32'sd424186, 32'sd325302,
32'sd469733, 32'sd757109, 32'sd599816, 32'sd115116, 32'sd162738, 32'sd247518, 32'sd519782, 32'sd289710, 32'sd35223, 32'sd7195,
32'sd115790, 32'sd137715, 32'sd401285, 32'sd81267, 32'sd96342, 32'sd339568, 32'sd706333, 32'sd10357, 32'sd449010, 32'sd63389,
32'sd133777, 32'sd123753, 32'sd153105, 32'sd136246, 32'sd509998, 32'sd285974, 32'sd98610, 32'sd102476, 32'sd132668, 32'sd190272,
32'sd680630, 32'sd221030, 32'sd237006, 32'sd187041, 32'sd278688, 32'sd159773, 32'sd265963, 32'sd391966, 32'sd1250517, 32'sd193230,
32'sd116989, 32'sd423512, 32'sd205055, 32'sd289851, 32'sd306649, 32'sd160799, 32'sd578155, 32'sd319419, 32'sd368154, 32'sd144759,
32'sd55205, 32'sd230548, 32'sd131558, 32'sd483522, 32'sd71115, 32'sd1263, 32'sd197828, 32'sd532933, 32'sd145687, 32'sd228048,
32'sd821857, 32'sd80565, 32'sd221852, 32'sd358650, 32'sd91134, 32'sd398406, 32'sd43054, 32'sd66579, 32'sd70560, 32'sd44590,
32'sd43295, 32'sd466203, 32'sd982509, 32'sd176090, 32'sd332552, 32'sd606631, 32'sd152720, 32'sd314700, 32'sd244757, 32'sd470739,
32'sd201502, 32'sd243686, 32'sd696373, 32'sd319105, 32'sd215911, 32'sd473082, 32'sd306823, 32'sd743980, 32'sd110999, 32'sd232929,
32'sd83570, 32'sd514, 32'sd610215, 32'sd429187, 32'sd460382, 32'sd154791, 32'sd160619, 32'sd5397, 32'sd768596, 32'sd762722,
32'sd137399, 32'sd20321, 32'sd36451, 32'sd279022, 32'sd2610, 32'sd841470, 32'sd562974, 32'sd23100, 32'sd24627, 32'sd329370,
32'sd886844, 32'sd50340, 32'sd220758, 32'sd257708, 32'sd246524, 32'sd142280, 32'sd335436, 32'sd161463, 32'sd127088, 32'sd2035,
32'sd116892, 32'sd619381, 32'sd132118, 32'sd356839, 32'sd927225, 32'sd321935, 32'sd23369, 32'sd479110, 32'sd80721, 32'sd194068,
32'sd146867, 32'sd5124, 32'sd97905, 32'sd692523, 32'sd389655, 32'sd692954, 32'sd668562, 32'sd255882, 32'sd375520, 32'sd501178,
32'sd122112, 32'sd655914, 32'sd29595, 32'sd303447, 32'sd630388, 32'sd192442, 32'sd99931, 32'sd382935, 32'sd766565, 32'sd282169,
32'sd364992, 32'sd479030, 32'sd110228, 32'sd222809, 32'sd53755, 32'sd531379, 32'sd83373, 32'sd1147146, 32'sd214999, 32'sd88012,
32'sd344141, 32'sd444942, 32'sd660482, 32'sd579087, 32'sd883286, 32'sd118758, 32'sd145554, 32'sd55572, 32'sd161305, 32'sd852323,
32'sd638224, 32'sd138029, 32'sd54566, 32'sd499877, 32'sd646234, 32'sd80056, 32'sd88323, 32'sd247917, 32'sd321837, 32'sd123402,
32'sd811927, 32'sd70279, 32'sd507867, 32'sd791042, 32'sd119210, 32'sd208419, 32'sd46056, 32'sd174601, 32'sd1241783, 32'sd34047,
32'sd498780, 32'sd351816, 32'sd133854, 32'sd39864, 32'sd697525, 32'sd497604, 32'sd310263, 32'sd97944, 32'sd213093, 32'sd72249,
32'sd22432, 32'sd181113, 32'sd367263, 32'sd287114, 32'sd211845, 32'sd136339, 32'sd690205, 32'sd786081, 32'sd557994, 32'sd12510,
32'sd94142, 32'sd222152, 32'sd153342, 32'sd170016, 32'sd1087290, 32'sd689212, 32'sd189718, 32'sd260254, 32'sd182748, 32'sd334790,
32'sd191156, 32'sd100908, 32'sd344199, 32'sd363276, 32'sd98001, 32'sd3591, 32'sd100519, 32'sd482970, 32'sd534301, 32'sd379127,
32'sd1012258, 32'sd295450, 32'sd350280, 32'sd168072, 32'sd70775, 32'sd587938, 32'sd567333, 32'sd56795, 32'sd29230, 32'sd398728,
32'sd266084, 32'sd123057, 32'sd90005, 32'sd756138, 32'sd732877, 32'sd261793, 32'sd9624, 32'sd681029, 32'sd196855, 32'sd718190,
32'sd303660, 32'sd96336, 32'sd226636, 32'sd299908, 32'sd141357, 32'sd259686, 32'sd35941, 32'sd305923, 32'sd28549, 32'sd338424,
32'sd1016118, 32'sd193903, 32'sd417120, 32'sd82192, 32'sd37529, 32'sd248836, 32'sd638454, 32'sd251030, 32'sd384434, 32'sd337240,
32'sd52610, 32'sd275759, 32'sd187645, 32'sd1038941, 32'sd14560, 32'sd455642, 32'sd40204, 32'sd1037089, 32'sd505045, 32'sd185765,
32'sd82070, 32'sd40457, 32'sd86006, 32'sd157717, 32'sd186541, 32'sd137709, 32'sd405072, 32'sd57944, 32'sd216000, 32'sd226778,
32'sd139207, 32'sd30158, 32'sd18644, 32'sd329055, 32'sd115443, 32'sd78118, 32'sd72674, 32'sd168290, 32'sd17278, 32'sd48090,
32'sd52006, 32'sd440569, 32'sd771249, 32'sd57015, 32'sd90560, 32'sd513017, 32'sd60061, 32'sd121769, 32'sd60377, 32'sd98118,
32'sd55532, 32'sd76761, 32'sd92960, 32'sd197609, 32'sd17471, 32'sd585647, 32'sd561856, 32'sd1105902, 32'sd356639, 32'sd236794,
32'sd120500, 32'sd255051, 32'sd301003, 32'sd34886, 32'sd94684, 32'sd96900, 32'sd20942, 32'sd295926, 32'sd157347, 32'sd668449,
32'sd686982, 32'sd44053, 32'sd445116, 32'sd226211, 32'sd405679, 32'sd27423, 32'sd492303, 32'sd439473, 32'sd136157, 32'sd123814,
32'sd156961, 32'sd136828, 32'sd366887, 32'sd388682, 32'sd413463, 32'sd817937, 32'sd352827, 32'sd460258, 32'sd96267, 32'sd88777,
32'sd468608, 32'sd88200, 32'sd468609, 32'sd619651, 32'sd5180, 32'sd643200, 32'sd976210, 32'sd9243, 32'sd76732, 32'sd622303,
32'sd535882, 32'sd98891, 32'sd385201, 32'sd282965, 32'sd546392, 32'sd257024, 32'sd12247, 32'sd783955, 32'sd369351, 32'sd712801,
32'sd113538, 32'sd78163, 32'sd470952, 32'sd314562, 32'sd60920, 32'sd250996, 32'sd246125, 32'sd294699, 32'sd111890, 32'sd108037,
32'sd84599, 32'sd558778, 32'sd67930, 32'sd313684, 32'sd52823, 32'sd128309, 32'sd153965, 32'sd174850, 32'sd199593, 32'sd179835,
32'sd748559, 32'sd85352, 32'sd346931, 32'sd474578, 32'sd525147, 32'sd134111, 32'sd256462, 32'sd815937, 32'sd149556, 32'sd167280,
32'sd132889, 32'sd473902, 32'sd169184, 32'sd261100, 32'sd110701, 32'sd123969, 32'sd77665, 32'sd310197, 32'sd45812, 32'sd160274,
32'sd226154, 32'sd584455, 32'sd573841, 32'sd141124, 32'sd38560, 32'sd930252, 32'sd666382, 32'sd268378, 32'sd233609, 32'sd841556,
32'sd147974, 32'sd163688, 32'sd387404, 32'sd154483, 32'sd489758, 32'sd21724, 32'sd55142, 32'sd112948, 32'sd429276, 32'sd317890,
32'sd137687, 32'sd1079132, 32'sd223456, 32'sd106664, 32'sd1086900, 32'sd66972, 32'sd26443, 32'sd25375, 32'sd160420, 32'sd64183,
32'sd148561, 32'sd94960, 32'sd58801, 32'sd6741, 32'sd496324, 32'sd481904, 32'sd73280, 32'sd99107, 32'sd648812, 32'sd747894,
32'sd110466, 32'sd614092, 32'sd341679, 32'sd266136, 32'sd144604, 32'sd356787, 32'sd241441, 32'sd616392, 32'sd801347, 32'sd298372,
32'sd515597, 32'sd30097, 32'sd117075, 32'sd127016, 32'sd630868, 32'sd8420, 32'sd100351, 32'sd280425, 32'sd156036, 32'sd748649,
32'sd60556, 32'sd32676, 32'sd397516, 32'sd207523, 32'sd275210, 32'sd208203, 32'sd891632, 32'sd136187, 32'sd126447, 32'sd125183,
32'sd625487, 32'sd425404, 32'sd143767, 32'sd281197, 32'sd341363, 32'sd167721, 32'sd70006, 32'sd402450, 32'sd127068, 32'sd67191,
32'sd335531, 32'sd313207, 32'sd857497, 32'sd27084, 32'sd119162, 32'sd82781, 32'sd406301, 32'sd107776, 32'sd25025, 32'sd26064,
32'sd381125, 32'sd151469, 32'sd420633, 32'sd271033, 32'sd29406, 32'sd811170, 32'sd320803, 32'sd99694, 32'sd293745, 32'sd533938,
32'sd286227, 32'sd320494, 32'sd1289087, 32'sd572578, 32'sd30069, 32'sd332535, 32'sd377892, 32'sd733523, 32'sd154992, 32'sd768701,
32'sd244560, 32'sd326713, 32'sd255810, 32'sd248746, 32'sd366361, 32'sd216631, 32'sd429016, 32'sd63067, 32'sd33433, 32'sd150362,
32'sd430845, 32'sd61831, 32'sd444669, 32'sd18986, 32'sd281549, 32'sd227518, 32'sd120541, 32'sd150999, 32'sd176140, 32'sd199303,
32'sd125793, 32'sd325722, 32'sd319791, 32'sd14919, 32'sd176878, 32'sd285433, 32'sd318269, 32'sd316524, 32'sd198358, 32'sd514693,
32'sd481653, 32'sd68030, 32'sd406067, 32'sd55950, 32'sd162694, 32'sd251974, 32'sd72090, 32'sd55730, 32'sd460257, 32'sd327110,
32'sd182301, 32'sd121669, 32'sd151172, 32'sd254054, 32'sd220409, 32'sd22230, 32'sd251369, 32'sd2300, 32'sd875178, 32'sd227641,
32'sd46326, 32'sd33740, 32'sd160038, 32'sd198320, 32'sd128677, 32'sd126111, 32'sd455939, 32'sd189720, 32'sd638237, 32'sd723948,
32'sd5564, 32'sd51178, 32'sd623312, 32'sd18462, 32'sd94306, 32'sd169872, 32'sd739290, 32'sd85155, 32'sd579982, 32'sd70168,
32'sd49088, 32'sd105433, 32'sd182429, 32'sd133917, 32'sd518350, 32'sd188910, 32'sd157379, 32'sd31585, 32'sd208534, 32'sd153519,
32'sd502214, 32'sd503325, 32'sd66499, 32'sd23653, 32'sd134232, 32'sd45196, 32'sd219249, 32'sd40367, 32'sd242895, 32'sd1021136,
32'sd294454, 32'sd944424, 32'sd53689, 32'sd435064, 32'sd103010, 32'sd20284, 32'sd331420, 32'sd28681, 32'sd558702, 32'sd342790,
32'sd464250, 32'sd469617, 32'sd13591, 32'sd1284536, 32'sd203241, 32'sd190826, 32'sd114666, 32'sd117099, 32'sd168614, 32'sd155167,
32'sd219503, 32'sd151488, 32'sd281991, 32'sd314761, 32'sd173514, 32'sd119891, 32'sd589610, 32'sd154072, 32'sd321426, 32'sd815652,
32'sd746146, 32'sd394063, 32'sd131610, 32'sd990822, 32'sd23707, 32'sd121184, 32'sd250480, 32'sd125721, 32'sd322300, 32'sd193592,
32'sd75842, 32'sd169302, 32'sd386440, 32'sd240574, 32'sd259423, 32'sd171223, 32'sd212101, 32'sd117036, 32'sd377625, 32'sd78734,
32'sd91086, 32'sd390395, 32'sd120743, 32'sd325602, 32'sd171713, 32'sd84478, 32'sd509518, 32'sd613392, 32'sd91325, 32'sd385974,
32'sd54759, 32'sd105617, 32'sd54733, 32'sd729138, 32'sd114203, 32'sd47490, 32'sd17656, 32'sd5776, 32'sd119324, 32'sd210168,
32'sd6839, 32'sd80626, 32'sd308719, 32'sd258597, 32'sd29132, 32'sd105196, 32'sd68332, 32'sd356295, 32'sd403823, 32'sd130149,
32'sd702502, 32'sd1081042, 32'sd177927, 32'sd949674, 32'sd173243, 32'sd40580, 32'sd22625, 32'sd345582, 32'sd198376, 32'sd524086,
32'sd46397, 32'sd341638, 32'sd1064063, 32'sd328126, 32'sd129162, 32'sd237017, 32'sd14840, 32'sd37145, 32'sd703442, 32'sd2604,
32'sd591868, 32'sd457699, 32'sd214596, 32'sd53558, 32'sd67755, 32'sd834254, 32'sd249910, 32'sd201348, 32'sd179654, 32'sd1039203,
32'sd792626, 32'sd68811, 32'sd23131, 32'sd265035, 32'sd171783, 32'sd27364, 32'sd225321, 32'sd145111, 32'sd305845, 32'sd716913,
32'sd576885, 32'sd434462, 32'sd12163, 32'sd108280, 32'sd8235, 32'sd357806, 32'sd218252, 32'sd187499, 32'sd257278, 32'sd81074,
32'sd252193, 32'sd89898, 32'sd264280, 32'sd722380, 32'sd150920, 32'sd125165, 32'sd66367, 32'sd228247, 32'sd392773, 32'sd67140,
32'sd549104, 32'sd5842, 32'sd102109, 32'sd162695, 32'sd45452, 32'sd702, 32'sd69718, 32'sd155295, 32'sd412428, 32'sd164528,
32'sd294614, 32'sd152991, 32'sd775151, 32'sd67265, 32'sd127947, 32'sd155728, 32'sd474151, 32'sd439704, 32'sd102318, 32'sd345521,
32'sd16127, 32'sd853694, 32'sd175940, 32'sd335921, 32'sd251713, 32'sd36974, 32'sd11649, 32'sd91303, 32'sd101561, 32'sd352711,
32'sd9533, 32'sd259734, 32'sd501876, 32'sd341557, 32'sd65042, 32'sd54673, 32'sd791058, 32'sd147266, 32'sd65959, 32'sd376621,
32'sd78762, 32'sd1166596, 32'sd741157, 32'sd321426, 32'sd326668, 32'sd67528, 32'sd97682, 32'sd288396, 32'sd287181, 32'sd70131,
32'sd221278, 32'sd21663, 32'sd398556, 32'sd162673, 32'sd638307, 32'sd329082, 32'sd310211, 32'sd212948

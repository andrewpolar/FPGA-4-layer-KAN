32'sd614147, 32'sd1148462, 32'sd768979, 32'sd1096568, 32'sd1091199, 32'sd579701, 32'sd692429, 32'sd639054, 32'sd976193, 32'sd514167, 32'sd688457, 32'sd1107619, 32'sd425348, 32'sd786385,
32'sd1122522, 32'sd477864, 32'sd746844, 32'sd615954, 32'sd1054512, 32'sd939147, 32'sd786877, 32'sd695560, 32'sd720639, 32'sd596423, 32'sd1195053, 32'sd604225, 32'sd735805, 32'sd1069637,
32'sd979535, 32'sd407956, 32'sd634228, 32'sd522910, 32'sd620882, 32'sd857334, 32'sd901577, 32'sd699382, 32'sd421163, 32'sd786312, 32'sd762446, 32'sd710645, 32'sd688761, 32'sd514551,
32'sd1156567, 32'sd577086, 32'sd1009881, 32'sd1174670, 32'sd563728, 32'sd845860, 32'sd436895, 32'sd559808, 32'sd1083024, 32'sd1075605, 32'sd854552, 32'sd767953, 32'sd685634, 32'sd954529
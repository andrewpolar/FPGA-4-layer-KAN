32'sd474262, 32'sd476106, 32'sd1032784, 32'sd598340, 32'sd448849, 32'sd1135210, 32'sd808148, 32'sd985912, 32'sd1123080, 32'sd520888, 32'sd880281, 32'sd638625, 32'sd944477, 32'sd973901,
32'sd870575, 32'sd691533, 32'sd710754, 32'sd825830, 32'sd1185392, 32'sd447912, 32'sd846475, 32'sd680724, 32'sd1188074, 32'sd1017571, 32'sd1158002, 32'sd636624, 32'sd617604, 32'sd738338,
32'sd1157661, 32'sd1108341, 32'sd935184, 32'sd818842, 32'sd432874, 32'sd1198186, 32'sd568913, 32'sd1144891, 32'sd805557, 32'sd469785, 32'sd1102149, 32'sd1074715, 32'sd583405, 32'sd1131718,
32'sd696445, 32'sd805141, 32'sd613558, 32'sd478339, 32'sd863073, 32'sd962383, 32'sd1199139, 32'sd534325, 32'sd812119, 32'sd496488, 32'sd423885, 32'sd954983, 32'sd840117, 32'sd975921,
32'sd526959, 32'sd570656, 32'sd424165, 32'sd847947, 32'sd459857, 32'sd538266, 32'sd1016607, 32'sd631685, 32'sd1199800, 32'sd413725, 32'sd885655, 32'sd976084, 32'sd885772, 32'sd815486,
32'sd936031, 32'sd738013, 32'sd479567, 32'sd600614, 32'sd407535, 32'sd790932, 32'sd593657, 32'sd464879, 32'sd528743, 32'sd1114396, 32'sd716024, 32'sd1007775, 32'sd416909, 32'sd508735,
32'sd870691, 32'sd939939, 32'sd1194470, 32'sd851328, 32'sd540052, 32'sd1013404, 32'sd903257, 32'sd527136, 32'sd636427, 32'sd1053783, 32'sd537039, 32'sd627658, 32'sd949576, 32'sd1172510,
32'sd1047668, 32'sd647290, 32'sd512578, 32'sd820819, 32'sd603672, 32'sd726269, 32'sd885695, 32'sd811458, 32'sd1204976, 32'sd414150, 32'sd703673, 32'sd533568, 32'sd524018, 32'sd1016004,
32'sd1116984, 32'sd785203, 32'sd1135767, 32'sd788672, 32'sd688297, 32'sd519208, 32'sd876753, 32'sd726544, 32'sd441936, 32'sd1022281, 32'sd888797, 32'sd475941, 32'sd418590, 32'sd1121219,
32'sd1066694, 32'sd441146, 32'sd449825, 32'sd1146188, 32'sd575828, 32'sd1180627, 32'sd743094, 32'sd886450, 32'sd458733, 32'sd630014, 32'sd1136589, 32'sd615441, 32'sd767584, 32'sd828322,
32'sd496792, 32'sd551744, 32'sd1047104, 32'sd739418, 32'sd865610, 32'sd734068, 32'sd903503, 32'sd1092537, 32'sd788762, 32'sd919597, 32'sd948994, 32'sd803905, 32'sd653419, 32'sd997321,
32'sd1144289, 32'sd977125, 32'sd1040275, 32'sd939914, 32'sd932255, 32'sd572674, 32'sd462243, 32'sd743107, 32'sd1097094, 32'sd1144603, 32'sd711027, 32'sd1116195, 32'sd748317, 32'sd476155,
32'sd1106443, 32'sd627530, 32'sd695033, 32'sd1072561, 32'sd609233, 32'sd874948, 32'sd973853, 32'sd897866, 32'sd674229, 32'sd508265, 32'sd934708, 32'sd541948, 32'sd488916, 32'sd692099,
32'sd635284, 32'sd813590, 32'sd1134519, 32'sd944056, 32'sd1035542, 32'sd1137220, 32'sd626829, 32'sd446900, 32'sd879208, 32'sd464268, 32'sd689603, 32'sd891195, 32'sd908943, 32'sd610047,
32'sd678611, 32'sd450781, 32'sd883056, 32'sd945175, 32'sd622041, 32'sd653842, 32'sd1200260, 32'sd501978, 32'sd828357, 32'sd925459, 32'sd915236, 32'sd679307, 32'sd541520, 32'sd521174,
32'sd456308, 32'sd493245, 32'sd1189044, 32'sd780047, 32'sd1136954, 32'sd454965, 32'sd807078, 32'sd902984, 32'sd801497, 32'sd877079, 32'sd837499, 32'sd738979, 32'sd501787, 32'sd726686,
32'sd460937, 32'sd554588, 32'sd740299, 32'sd581570, 32'sd805514, 32'sd771677, 32'sd422597, 32'sd1043730, 32'sd564401, 32'sd1105126, 32'sd954981, 32'sd1144939, 32'sd711949, 32'sd456617,
32'sd417415, 32'sd1010404, 32'sd745787, 32'sd621939, 32'sd734243, 32'sd780981, 32'sd424408, 32'sd781808, 32'sd977466, 32'sd558316, 32'sd414482, 32'sd508347, 32'sd430698, 32'sd1056442,
32'sd876114, 32'sd951831, 32'sd1136080, 32'sd413348, 32'sd664903, 32'sd1187452, 32'sd498673, 32'sd1058943, 32'sd877576, 32'sd594634, 32'sd641685, 32'sd689922, 32'sd767960, 32'sd723287,
32'sd483978, 32'sd513755, 32'sd671169, 32'sd1143351, 32'sd803154, 32'sd1076468, 32'sd854967, 32'sd960046, 32'sd1177060, 32'sd966431, 32'sd986315, 32'sd1062824, 32'sd526019, 32'sd533820,
32'sd1011152, 32'sd410146, 32'sd1104686, 32'sd661924, 32'sd463380, 32'sd774554, 32'sd721368, 32'sd489398, 32'sd647822, 32'sd1101324, 32'sd716594, 32'sd1171069, 32'sd923691, 32'sd953463,
32'sd403832, 32'sd642308, 32'sd414028, 32'sd717953, 32'sd843185, 32'sd964024, 32'sd1159511, 32'sd788973, 32'sd677494, 32'sd923720, 32'sd940356, 32'sd961514, 32'sd1081205, 32'sd1028787,
32'sd956056, 32'sd1140789, 32'sd617571, 32'sd952582, 32'sd865518, 32'sd977131, 32'sd925495, 32'sd502256, 32'sd639674, 32'sd1152278, 32'sd959558, 32'sd986459, 32'sd464972, 32'sd1019251,
32'sd552500, 32'sd999801, 32'sd900906, 32'sd892864, 32'sd802558, 32'sd810180, 32'sd663732, 32'sd1021951, 32'sd704816, 32'sd777853, 32'sd485210, 32'sd965289, 32'sd694627, 32'sd996082,
32'sd1186763, 32'sd1003710, 32'sd1168444, 32'sd1125179, 32'sd1069290, 32'sd784041, 32'sd510559, 32'sd831783, 32'sd784762, 32'sd424560, 32'sd892718, 32'sd1011923, 32'sd707835, 32'sd638333,
32'sd1150598, 32'sd1173352, 32'sd1104336, 32'sd1009707, 32'sd1103576, 32'sd1084650, 32'sd442937, 32'sd623581, 32'sd1053614, 32'sd481258, 32'sd1084106, 32'sd1125383, 32'sd802955, 32'sd1049145,
32'sd498862, 32'sd1016510, 32'sd1162756, 32'sd1147471, 32'sd1068157, 32'sd1023058, 32'sd957383, 32'sd1001135, 32'sd965202, 32'sd476601, 32'sd1151188, 32'sd740517, 32'sd901668, 32'sd499602,
32'sd984817, 32'sd919319, 32'sd1092700, 32'sd951199, 32'sd742956, 32'sd729607, 32'sd950608, 32'sd444696, 32'sd852703, 32'sd978498, 32'sd739492, 32'sd988536, 32'sd1067481, 32'sd1162190,
32'sd633687, 32'sd1009275, 32'sd942061, 32'sd737072, 32'sd730443, 32'sd1010104, 32'sd1153884, 32'sd886119, 32'sd1048449, 32'sd922671, 32'sd1139196, 32'sd738586, 32'sd494235, 32'sd1076948,
32'sd616129, 32'sd868307, 32'sd412016, 32'sd919493, 32'sd539717, 32'sd415581, 32'sd1030757, 32'sd858672, 32'sd524744, 32'sd775425, 32'sd1195136, 32'sd415172, 32'sd607764, 32'sd873862,
32'sd748553, 32'sd946020, 32'sd614849, 32'sd708821, 32'sd1085645, 32'sd601680, 32'sd958432, 32'sd410747, 32'sd514038, 32'sd626545, 32'sd1163269, 32'sd562549, 32'sd773373, 32'sd1071714,
32'sd830852, 32'sd635325, 32'sd643235, 32'sd705438, 32'sd947583, 32'sd696078, 32'sd1051473, 32'sd584888, 32'sd584592, 32'sd766269, 32'sd672829, 32'sd902752, 32'sd592247, 32'sd961395,
32'sd1164668, 32'sd409352, 32'sd972476, 32'sd759098, 32'sd602701, 32'sd670853, 32'sd801379, 32'sd1078495, 32'sd700546, 32'sd552194, 32'sd723508, 32'sd642385, 32'sd489606, 32'sd464320,
32'sd1082452, 32'sd976988, 32'sd1019664, 32'sd452470, 32'sd601581, 32'sd627519, 32'sd1035265, 32'sd428870, 32'sd1030265, 32'sd769125, 32'sd1069541, 32'sd677051, 32'sd972948, 32'sd436787,
32'sd901216, 32'sd478901, 32'sd788744, 32'sd514670, 32'sd487363, 32'sd735980, 32'sd516674, 32'sd1069431, 32'sd622042, 32'sd1010220, 32'sd1034777, 32'sd476653, 32'sd449278, 32'sd889608,
32'sd423764, 32'sd651986, 32'sd968858, 32'sd673961, 32'sd721688, 32'sd820316, 32'sd815523, 32'sd953588, 32'sd861857, 32'sd1131441, 32'sd1148922, 32'sd1004390, 32'sd778467, 32'sd887545,
32'sd806689, 32'sd1149616, 32'sd892121, 32'sd1158225, 32'sd469463, 32'sd915948, 32'sd1026526, 32'sd508931, 32'sd932185, 32'sd965959, 32'sd1164986, 32'sd863330, 32'sd1022142, 32'sd567915,
32'sd764213, 32'sd472138, 32'sd977192, 32'sd900133, 32'sd1021524, 32'sd630503, 32'sd674292, 32'sd611741, 32'sd1109301, 32'sd907823, 32'sd986863, 32'sd1005608, 32'sd469756, 32'sd932255,
32'sd688106, 32'sd1078879, 32'sd570023, 32'sd690778, 32'sd736759, 32'sd953787, 32'sd1070017, 32'sd1115801, 32'sd746736, 32'sd732685, 32'sd755051, 32'sd611384, 32'sd655847, 32'sd881128,
32'sd1011427, 32'sd869882, 32'sd1040098, 32'sd990774, 32'sd927480, 32'sd1019076, 32'sd803466, 32'sd805968, 32'sd974208, 32'sd561163, 32'sd827413, 32'sd411442, 32'sd917127, 32'sd430715,
32'sd1195894, 32'sd1013653, 32'sd627654, 32'sd1168383, 32'sd692870, 32'sd754024, 32'sd516566, 32'sd925446, 32'sd994051, 32'sd1197373, 32'sd919997, 32'sd443262, 32'sd597084, 32'sd1163260,
32'sd450109, 32'sd832027, 32'sd1048383, 32'sd515611, 32'sd1136989, 32'sd590226, 32'sd1058702, 32'sd844759, 32'sd793756, 32'sd522059, 32'sd535590, 32'sd1122073, 32'sd1053687, 32'sd1072561,
32'sd1010136, 32'sd568308, 32'sd1067384, 32'sd1143321, 32'sd897043, 32'sd1049897, 32'sd1127945, 32'sd451238, 32'sd1065385, 32'sd1007649, 32'sd602821, 32'sd807102, 32'sd941006, 32'sd1133339,
32'sd1047246, 32'sd975336, 32'sd456287, 32'sd1105067, 32'sd726550, 32'sd707473, 32'sd644751, 32'sd655030, 32'sd999436, 32'sd679975, 32'sd465863, 32'sd1123067, 32'sd1091678, 32'sd1081191